magic
tech scmos
timestamp 1714289837
<< metal1 >>
rect -1476 3377 -1472 3381
rect -1389 3377 -1385 3392
rect -1476 3373 -1385 3377
rect -1176 3374 -1172 3380
rect -1089 3374 -1085 3392
rect -1176 3370 -1085 3374
rect -876 3374 -872 3380
rect -789 3374 -785 3392
rect -876 3370 -785 3374
rect -576 3374 -572 3379
rect -489 3374 -485 3392
rect -576 3370 -485 3374
rect -276 3371 -272 3380
rect -189 3371 -185 3392
rect -276 3367 -185 3371
rect 25 3374 29 3380
rect 111 3374 115 3392
rect 25 3370 115 3374
rect 435 2619 458 3407
rect 924 3377 928 3380
rect 1011 3377 1015 3392
rect 924 3373 1015 3377
rect 1224 3376 1228 3381
rect 1311 3376 1315 3392
rect 1224 3372 1315 3376
rect 1524 3375 1528 3380
rect 1611 3375 1615 3392
rect 1524 3371 1615 3375
rect 1824 3373 1828 3379
rect 1911 3373 1915 3392
rect 1824 3369 1915 3373
rect 2123 3366 2127 3380
rect 2211 3366 2215 3393
rect 2123 3362 2215 3366
rect 798 3330 799 3336
rect 805 3330 829 3336
rect 799 3315 800 3320
rect 805 3315 812 3320
rect 784 3296 789 3300
rect 763 3282 774 3283
rect 769 3276 774 3282
rect 749 3261 756 3266
rect 729 3245 738 3246
rect 734 3240 738 3245
rect 733 3143 738 3240
rect 751 3155 756 3261
rect 768 3173 774 3276
rect 785 3186 789 3296
rect 807 3205 812 3315
rect 823 3223 829 3330
rect 823 3217 1450 3223
rect 807 3202 1622 3205
rect 807 3200 1617 3202
rect 1621 3197 1622 3202
rect 785 3182 1786 3186
rect 768 3167 1954 3173
rect 751 3150 2058 3155
rect 733 3138 2162 3143
rect 435 2596 585 2619
rect 2535 2604 2558 3407
rect 2727 3378 2729 3383
rect 2725 3376 2729 3378
rect 2811 3376 2815 3392
rect 2725 3372 2815 3376
rect 3025 3374 3029 3379
rect 3111 3374 3115 3392
rect 3025 3370 3115 3374
rect 3266 3211 3292 3215
rect 3266 3129 3270 3211
rect 3266 3125 3281 3129
rect 3266 2911 3292 2915
rect 3266 2828 3270 2911
rect 3266 2824 3280 2828
rect 562 2528 585 2596
rect 2384 2581 2558 2604
rect 3267 2611 3292 2615
rect 2384 2529 2407 2581
rect 3267 2529 3271 2611
rect 3267 2525 3282 2529
rect 3259 2311 3292 2315
rect 3259 2229 3263 2311
rect 3259 2225 3281 2229
rect -624 2096 -557 2109
rect -624 2053 -611 2096
rect -1502 2040 -611 2053
rect 3263 2011 3292 2015
rect 3263 1928 3267 2011
rect 3263 1924 3282 1928
rect 2441 1746 3302 1759
rect -1492 1411 -1461 1415
rect -1465 1328 -1461 1411
rect -1480 1324 -1461 1328
rect 3269 1411 3293 1415
rect 3269 1329 3273 1411
rect 3269 1325 3282 1329
rect -1494 1111 -1464 1115
rect -1468 1030 -1464 1111
rect -1480 1026 -1464 1030
rect 3269 1111 3292 1115
rect 3269 1029 3273 1111
rect 3269 1025 3280 1029
rect -1492 811 -1460 815
rect -1464 729 -1460 811
rect -1483 725 -1460 729
rect 3268 811 3292 815
rect 3268 729 3272 811
rect 3268 725 3279 729
rect -1492 511 -1464 515
rect -1468 428 -1464 511
rect -1480 424 -1464 428
rect 3266 511 3292 515
rect 3266 429 3270 511
rect 3266 425 3281 429
rect -1502 246 -556 259
rect 3264 211 3292 215
rect 3264 129 3268 211
rect 3264 125 3281 129
rect -1480 72 -1468 76
rect -1472 -11 -1468 72
rect -1492 -15 -1468 -11
rect 2511 -54 3302 -41
rect 2511 -70 2524 -54
rect 2439 -83 2524 -70
rect -1495 -389 -1466 -385
rect -1470 -471 -1466 -389
rect 3268 -389 3292 -385
rect -1480 -475 -1466 -471
rect -188 -510 -165 -464
rect -188 -533 -142 -510
rect 1717 -522 1740 -466
rect 3268 -471 3272 -389
rect 3268 -475 3281 -471
rect -1493 -689 -1466 -685
rect -1488 -776 -1487 -772
rect -1470 -772 -1466 -689
rect -1481 -776 -1466 -772
rect -1492 -989 -1467 -985
rect -1471 -1072 -1467 -989
rect -1480 -1076 -1467 -1072
rect -1492 -1289 -1454 -1285
rect -1458 -1359 -1454 -1289
rect -1175 -1372 -1085 -1368
rect -1175 -1380 -1171 -1372
rect -1089 -1392 -1085 -1372
rect -875 -1373 -785 -1369
rect -875 -1381 -871 -1373
rect -789 -1392 -785 -1373
rect -576 -1375 -485 -1371
rect -576 -1380 -572 -1375
rect -489 -1392 -485 -1375
rect -165 -1407 -142 -533
rect 1635 -545 1740 -522
rect 24 -1368 115 -1364
rect 24 -1379 28 -1368
rect 111 -1392 115 -1368
rect 325 -1374 415 -1370
rect 924 -1371 1015 -1367
rect 325 -1380 329 -1374
rect 411 -1392 415 -1374
rect 624 -1376 715 -1372
rect 624 -1382 628 -1376
rect 711 -1393 715 -1376
rect 924 -1385 928 -1371
rect 1011 -1392 1015 -1371
rect 1225 -1370 1315 -1366
rect 1225 -1379 1229 -1370
rect 1311 -1392 1315 -1370
rect 1635 -1407 1658 -545
rect 3261 -689 3292 -685
rect 3261 -772 3265 -689
rect 3261 -776 3281 -772
rect 3267 -989 3292 -985
rect 3267 -1073 3271 -989
rect 3267 -1077 3280 -1073
rect 3273 -1289 3292 -1285
rect 2424 -1370 2515 -1366
rect 1824 -1375 1915 -1371
rect 1824 -1383 1828 -1375
rect 1911 -1392 1915 -1375
rect 2124 -1375 2215 -1371
rect 2124 -1380 2128 -1375
rect 2211 -1392 2215 -1375
rect 2424 -1380 2428 -1370
rect 2511 -1392 2515 -1370
rect 2725 -1373 2815 -1369
rect 3273 -1371 3277 -1289
rect 2725 -1381 2729 -1373
rect 2811 -1392 2815 -1373
rect 3024 -1377 3115 -1373
rect 3273 -1375 3280 -1371
rect 3024 -1381 3028 -1377
rect 3111 -1392 3115 -1377
<< m2contact >>
rect -1477 3381 -1471 3387
rect -1177 3380 -1171 3386
rect -877 3380 -871 3386
rect -577 3379 -571 3385
rect -277 3380 -271 3386
rect 24 3380 30 3386
rect 923 3380 929 3385
rect 1222 3381 1229 3386
rect 1523 3380 1529 3386
rect 1823 3379 1829 3385
rect 2122 3380 2128 3386
rect 799 3330 805 3336
rect 800 3315 805 3320
rect 780 3296 784 3300
rect 763 3276 769 3282
rect 744 3261 749 3266
rect 729 3240 734 3245
rect 1450 3217 1454 3223
rect 1617 3197 1621 3202
rect 1786 3182 1790 3186
rect 1954 3167 1958 3173
rect 2058 3150 2062 3155
rect 2162 3138 2166 3143
rect 2721 3378 2727 3384
rect 3024 3379 3030 3385
rect 3281 3124 3287 3130
rect 3280 2823 3286 2829
rect 3282 2524 3288 2530
rect 3281 2224 3287 2230
rect -557 2093 -537 2113
rect 3282 1923 3288 1929
rect 2421 1743 2441 1763
rect -1486 1323 -1480 1329
rect 3282 1324 3288 1330
rect -1486 1025 -1480 1031
rect 3280 1024 3286 1030
rect -1489 724 -1483 730
rect 3279 724 3285 730
rect -1486 423 -1480 429
rect 3281 424 3287 430
rect -556 243 -536 263
rect 3281 124 3287 130
rect -1486 71 -1480 77
rect 2419 -86 2439 -66
rect -1486 -476 -1480 -470
rect 3281 -476 3287 -470
rect -1487 -777 -1481 -771
rect -1486 -1077 -1480 -1071
rect -1459 -1365 -1453 -1359
rect -1176 -1386 -1170 -1380
rect -876 -1387 -870 -1381
rect -577 -1386 -571 -1380
rect 23 -1385 29 -1379
rect 324 -1386 330 -1380
rect 623 -1388 629 -1382
rect 1224 -1385 1230 -1379
rect 3281 -777 3287 -771
rect 3280 -1078 3286 -1072
rect 1823 -1389 1829 -1383
rect 2123 -1386 2129 -1380
rect 2423 -1386 2429 -1380
rect 2723 -1387 2729 -1381
rect 3280 -1376 3286 -1370
rect 3023 -1387 3029 -1381
<< metal2 >>
rect -1484 3359 -1465 3362
rect -1468 3345 -1465 3359
rect -1451 3355 -1448 3383
rect -1451 3352 -1201 3355
rect -1468 3342 -1293 3345
rect -1492 3194 -1465 3200
rect -1471 3129 -1465 3194
rect -1488 3123 -1465 3129
rect -1485 3058 -1302 3061
rect -1492 2894 -1468 2900
rect -1474 2829 -1468 2894
rect -1487 2823 -1468 2829
rect -1484 2758 -1312 2761
rect -1491 2594 -1461 2600
rect -1467 2529 -1461 2594
rect -1487 2523 -1461 2529
rect -1484 2457 -1325 2460
rect -1492 2294 -1466 2300
rect -1472 2229 -1466 2294
rect -1487 2223 -1466 2229
rect -1487 1871 -1456 1877
rect -1462 1805 -1456 1871
rect -1492 1799 -1456 1805
rect -1486 1634 -1336 1637
rect -1484 1345 -1347 1348
rect -1487 1044 -1360 1047
rect -1484 744 -1373 747
rect -1485 445 -1385 448
rect -1486 49 -1397 52
rect -1486 -454 -1414 -451
rect -1488 -754 -1430 -751
rect -1486 -1052 -1444 -1049
rect -1447 -1258 -1444 -1052
rect -1433 -1242 -1430 -754
rect -1417 -1233 -1414 -454
rect -1400 -1222 -1397 49
rect -1388 -1213 -1385 445
rect -1376 -1205 -1373 744
rect -1363 -1197 -1360 1044
rect -1350 -1188 -1347 1345
rect -1339 -1177 -1336 1634
rect -1328 583 -1325 2457
rect -1315 643 -1312 2758
rect -1305 963 -1302 3058
rect -1296 1703 -1293 3342
rect -1204 3244 -1201 3352
rect -1152 3264 -1149 3384
rect -854 3281 -850 3385
rect -552 3299 -549 3385
rect -253 3319 -249 3384
rect 44 3335 49 3384
rect 623 3377 629 3387
rect 694 3377 700 3392
rect 623 3371 700 3377
rect 44 3330 799 3335
rect -253 3315 800 3319
rect -552 3296 780 3299
rect -854 3277 763 3281
rect -1152 3261 744 3264
rect -1204 3241 729 3244
rect 860 3159 863 3386
rect 946 3370 949 3384
rect 946 3367 1046 3370
rect 860 3156 990 3159
rect 987 2545 990 3156
rect 1043 2545 1046 3367
rect 1247 3362 1250 3385
rect 1059 3359 1250 3362
rect 1059 2545 1062 3359
rect 1547 3341 1550 3384
rect 1075 3338 1550 3341
rect 1075 2545 1078 3338
rect 1848 3313 1851 3383
rect 1163 3310 1851 3313
rect 1163 2545 1166 3310
rect 2148 3297 2151 3385
rect 1179 3294 2151 3297
rect 1179 2545 1182 3294
rect 2747 3278 2750 3385
rect 1203 3275 2750 3278
rect 1203 2545 1206 3275
rect 3045 3259 3048 3384
rect 1371 3256 3048 3259
rect 1371 2545 1374 3256
rect 2267 3236 3260 3239
rect 1451 2545 1454 3217
rect 1621 3197 1622 3202
rect 1619 2545 1622 3197
rect 1787 2545 1790 3182
rect 1955 2545 1958 3167
rect 2059 2545 2062 3150
rect 2163 2545 2166 3138
rect 2267 2545 2270 3236
rect 3257 3150 3260 3236
rect 3257 3147 3285 3150
rect 3063 2847 3286 2852
rect 3063 1855 3068 2847
rect 2519 1850 3068 1855
rect 3080 2546 3286 2551
rect 2521 1720 2523 1724
rect 3080 1724 3085 2546
rect 2528 1720 3085 1724
rect 2521 1719 3085 1720
rect 3094 2252 3274 2257
rect -1296 1700 -626 1703
rect 3094 1615 3099 2252
rect 3269 2251 3274 2252
rect 3269 2246 3284 2251
rect 2516 1610 3099 1615
rect 3114 1947 3286 1951
rect 3114 1524 3118 1947
rect 2523 1520 3118 1524
rect 3255 1345 3286 1349
rect 3255 1344 3259 1345
rect 2506 1340 3259 1344
rect 2507 1210 3259 1213
rect 2518 1070 3241 1073
rect -1305 960 -641 963
rect 3238 751 3241 1070
rect 3256 1051 3259 1210
rect 3256 1048 3284 1051
rect 3238 748 3285 751
rect 2522 650 3240 654
rect -1315 640 -645 643
rect 2530 610 3222 614
rect 2534 590 2535 594
rect 2540 590 3202 594
rect -1328 580 -632 583
rect -627 580 -626 583
rect 898 548 2467 568
rect 2540 540 2541 544
rect 2546 540 3184 544
rect 2556 520 3169 524
rect 2557 500 3157 503
rect 2532 -280 2534 -277
rect 2539 -280 3130 -277
rect 2543 -370 2544 -366
rect 2549 -370 2731 -366
rect -261 -1177 -258 -489
rect -1339 -1180 -258 -1177
rect 283 -1188 286 -489
rect -1350 -1191 286 -1188
rect 379 -1197 382 -489
rect -1363 -1200 382 -1197
rect 395 -1205 398 -489
rect -1376 -1208 398 -1205
rect 411 -1213 414 -489
rect -1388 -1216 414 -1213
rect 435 -1222 438 -489
rect -1400 -1225 438 -1222
rect 539 -1233 542 -489
rect -1417 -1236 542 -1233
rect 555 -1242 558 -489
rect -1433 -1245 558 -1242
rect 731 -1258 734 -489
rect -1447 -1261 734 -1258
rect 907 -1270 910 -489
rect -1468 -1273 910 -1270
rect -1468 -1348 -1465 -1273
rect 971 -1278 974 -489
rect -1483 -1351 -1465 -1348
rect -1238 -1281 974 -1278
rect -1487 -1365 -1459 -1359
rect -1487 -1377 -1481 -1365
rect -1469 -1375 -1399 -1369
rect -1469 -1381 -1463 -1375
rect -1477 -1387 -1463 -1381
rect -1405 -1390 -1399 -1375
rect -1238 -1384 -1235 -1281
rect 1067 -1287 1070 -489
rect -1154 -1290 1070 -1287
rect -1154 -1385 -1151 -1290
rect 1083 -1296 1086 -489
rect -851 -1299 1086 -1296
rect -851 -1386 -848 -1299
rect 1115 -1305 1118 -489
rect -552 -1308 1118 -1305
rect -552 -1384 -549 -1308
rect 1219 -1313 1222 -489
rect 47 -1316 1222 -1313
rect 47 -1387 50 -1316
rect 1235 -1321 1238 -489
rect 346 -1324 1238 -1321
rect 346 -1388 349 -1324
rect 1379 -1330 1382 -489
rect 649 -1333 1382 -1330
rect 649 -1382 652 -1333
rect 1619 -1340 1622 -489
rect 945 -1343 1622 -1340
rect 945 -1384 948 -1343
rect 1787 -1354 1790 -489
rect 1245 -1357 1790 -1354
rect 1245 -1384 1248 -1357
rect 1963 -1366 1966 -489
rect 2107 -1339 2110 -489
rect 2243 -1320 2246 -489
rect 2727 -1228 2731 -370
rect 2727 -1232 2751 -1228
rect 2243 -1323 2452 -1320
rect 2107 -1342 2154 -1339
rect 1847 -1369 1966 -1366
rect 1847 -1386 1850 -1369
rect 2151 -1376 2154 -1342
rect 2144 -1383 2154 -1376
rect 2144 -1390 2153 -1383
rect 2449 -1386 2452 -1323
rect 2747 -1385 2751 -1232
rect 3127 -1366 3130 -280
rect 3154 -1076 3157 500
rect 3165 -1047 3169 520
rect 3180 -745 3184 540
rect 3198 -446 3202 590
rect 3218 153 3222 610
rect 3236 451 3240 650
rect 3236 447 3284 451
rect 3218 149 3287 153
rect 3198 -450 3275 -446
rect 3271 -454 3286 -450
rect 3180 -749 3285 -745
rect 3165 -1051 3287 -1047
rect 3154 -1079 3254 -1076
rect 3251 -1349 3254 -1079
rect 3251 -1352 3282 -1349
rect 3047 -1369 3130 -1366
rect 3047 -1385 3050 -1369
<< m3contact >>
rect 2514 1850 2519 1855
rect 2523 1720 2528 1725
rect -626 1700 -621 1705
rect 2511 1610 2516 1615
rect 2518 1520 2523 1525
rect 2501 1340 2506 1345
rect 2502 1210 2507 1215
rect 2513 1070 2518 1075
rect -641 960 -636 965
rect 2517 650 2522 655
rect -645 640 -640 645
rect 2525 610 2530 615
rect 2535 590 2540 595
rect -632 580 -627 585
rect 2541 540 2546 545
rect 2551 520 2556 525
rect 2552 500 2557 505
rect 2534 -280 2539 -275
rect 2544 -370 2549 -365
<< metal3 >>
rect 2513 1855 2520 1856
rect 2476 1850 2514 1855
rect 2519 1850 2520 1855
rect 2513 1849 2520 1850
rect 2522 1725 2529 1726
rect 2476 1720 2523 1725
rect 2528 1720 2529 1725
rect 2522 1719 2529 1720
rect -627 1705 -620 1706
rect -627 1700 -626 1705
rect -621 1700 -594 1705
rect -627 1699 -620 1700
rect 2510 1615 2517 1616
rect 2475 1610 2511 1615
rect 2516 1610 2517 1615
rect 2510 1609 2517 1610
rect 2517 1525 2524 1526
rect 2476 1520 2518 1525
rect 2523 1520 2524 1525
rect 2517 1519 2524 1520
rect 2500 1345 2507 1346
rect 2476 1340 2501 1345
rect 2506 1340 2507 1345
rect 2500 1339 2507 1340
rect 2501 1215 2508 1216
rect 2476 1210 2502 1215
rect 2507 1210 2508 1215
rect 2501 1209 2508 1210
rect 2512 1075 2519 1076
rect 2476 1070 2513 1075
rect 2518 1070 2519 1075
rect 2512 1069 2519 1070
rect -642 965 -635 966
rect -642 960 -641 965
rect -636 960 -594 965
rect -642 959 -635 960
rect 2516 655 2523 656
rect 2476 650 2517 655
rect 2522 650 2523 655
rect 2516 649 2523 650
rect -646 645 -639 646
rect -646 640 -645 645
rect -640 640 -594 645
rect -646 639 -639 640
rect 2524 615 2531 616
rect 2476 610 2525 615
rect 2530 610 2531 615
rect 2524 609 2531 610
rect 2534 595 2541 596
rect 2476 590 2535 595
rect 2540 590 2541 595
rect 2534 589 2541 590
rect -633 585 -626 586
rect -633 580 -632 585
rect -627 580 -594 585
rect -633 579 -626 580
rect 2540 545 2547 546
rect 2476 540 2541 545
rect 2546 540 2547 545
rect 2540 539 2547 540
rect 2550 525 2557 526
rect 2476 520 2551 525
rect 2556 520 2557 525
rect 2550 519 2557 520
rect 2551 505 2558 506
rect 2476 500 2552 505
rect 2557 500 2558 505
rect 2551 499 2558 500
rect 2533 -275 2540 -274
rect 2476 -280 2534 -275
rect 2539 -280 2540 -275
rect 2533 -281 2540 -280
rect 2543 -365 2550 -364
rect 2476 -370 2544 -365
rect 2549 -370 2550 -365
rect 2543 -371 2550 -370
use PadFC  16_0
timestamp 1681001061
transform 1 0 -2500 0 1 3400
box 327 -3 1003 673
use PadFC  16_1
timestamp 1681001061
transform 0 1 3300 -1 0 4400
box 327 -3 1003 673
use PadFC  16_2
timestamp 1681001061
transform 0 -1 -1500 1 0 -2400
box 327 -3 1003 673
use PadFC  16_3
timestamp 1681001061
transform -1 0 4300 0 -1 -1400
box 327 -3 1003 673
use PadBiDir  17_0
timestamp 1711830429
transform 1 0 -1500 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_1
timestamp 1711830429
transform 1 0 -1200 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_2
timestamp 1711830429
transform 1 0 -900 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_3
timestamp 1711830429
transform 1 0 -600 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_4
timestamp 1711830429
transform 1 0 -300 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_5
timestamp 1711830429
transform 1 0 0 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_6
timestamp 1711830429
transform 1 0 600 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_7
timestamp 1711830429
transform 1 0 900 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_8
timestamp 1711830429
transform 1 0 1200 0 1 3400
box -36 -19 303 1000
use PadBiDir  17_9
timestamp 1711830429
transform 0 -1 -1500 1 0 3100
box -36 -19 303 1000
use PadBiDir  17_10
timestamp 1711830429
transform 0 -1 -1500 1 0 2800
box -36 -19 303 1000
use PadBiDir  17_11
timestamp 1711830429
transform 0 -1 -1500 1 0 2500
box -36 -19 303 1000
use PadBiDir  17_12
timestamp 1711830429
transform 0 -1 -1500 1 0 2200
box -36 -19 303 1000
use PadBiDir  17_13
timestamp 1711830429
transform 0 -1 -1500 -1 0 1900
box -36 -19 303 1000
use PadBiDir  17_14
timestamp 1711830429
transform 0 -1 -1500 1 0 -500
box -36 -19 303 1000
use PadBiDir  17_15
timestamp 1711830429
transform 0 -1 -1500 1 0 -800
box -36 -19 303 1000
use PadBiDir  17_16
timestamp 1711830429
transform 0 -1 -1500 1 0 -1100
box -36 -19 303 1000
use PadBiDir  17_17
timestamp 1711830429
transform 0 1 3300 1 0 3100
box -36 -19 303 1000
use PadBiDir  17_18
timestamp 1711830429
transform 0 1 3300 1 0 2800
box -36 -19 303 1000
use PadBiDir  17_19
timestamp 1711830429
transform 0 1 3300 1 0 2500
box -36 -19 303 1000
use PadBiDir  17_20
timestamp 1711830429
transform 0 1 3300 1 0 2200
box -36 -19 303 1000
use PadBiDir  17_21
timestamp 1711830429
transform 0 1 3300 1 0 1900
box -36 -19 303 1000
use PadBiDir  17_22
timestamp 1711830429
transform 0 1 3300 1 0 -500
box -36 -19 303 1000
use PadBiDir  17_23
timestamp 1711830429
transform 0 1 3300 1 0 -800
box -36 -19 303 1000
use PadBiDir  17_24
timestamp 1711830429
transform 0 1 3300 1 0 -1100
box -36 -19 303 1000
use PadBiDir  17_25
timestamp 1711830429
transform 0 -1 -1500 1 0 -1400
box -36 -19 303 1000
use PadBiDir  17_26
timestamp 1711830429
transform 1 0 -1500 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_27
timestamp 1711830429
transform 1 0 -1200 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_28
timestamp 1711830429
transform 1 0 -900 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_29
timestamp 1711830429
transform 1 0 -600 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_30
timestamp 1711830429
transform 1 0 0 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_31
timestamp 1711830429
transform 1 0 300 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_32
timestamp 1711830429
transform 1 0 600 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_33
timestamp 1711830429
transform 1 0 900 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  17_34
timestamp 1711830429
transform 0 1 3300 1 0 -1400
box -36 -19 303 1000
use PadBiDir  17_35
timestamp 1711830429
transform 1 0 1200 0 -1 -1400
box -36 -19 303 1000
use PadVdd  18_0
timestamp 1711831643
transform 1 0 300 0 1 3400
box -3 -16 303 1000
use PadVdd  18_1
timestamp 1711831643
transform 1 0 -300 0 -1 -1400
box -3 -16 303 1000
use PadGnd  19_0
timestamp 1711831454
transform 0 -1 -1500 -1 0 2200
box -3 -11 303 1000
use PadGnd  19_1
timestamp 1711831454
transform 0 1 3300 -1 0 1900
box -3 -11 303 1000
use PadBiDir  PadBiDir_0
timestamp 1711830429
transform 1 0 1500 0 1 3400
box -36 -19 303 1000
use PadBiDir  PadBiDir_1
timestamp 1711830429
transform 1 0 1800 0 1 3400
box -36 -19 303 1000
use PadBiDir  PadBiDir_2
timestamp 1711830429
transform 1 0 2100 0 1 3400
box -36 -19 303 1000
use PadBiDir  PadBiDir_3
timestamp 1711830429
transform 1 0 2700 0 1 3400
box -36 -19 303 1000
use PadBiDir  PadBiDir_4
timestamp 1711830429
transform 1 0 3000 0 1 3400
box -36 -19 303 1000
use PadBiDir  PadBiDir_5
timestamp 1711830429
transform 1 0 1800 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  PadBiDir_6
timestamp 1711830429
transform 1 0 2100 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  PadBiDir_7
timestamp 1711830429
transform 1 0 2400 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  PadBiDir_8
timestamp 1711830429
transform 1 0 2700 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  PadBiDir_9
timestamp 1711830429
transform 1 0 3000 0 -1 -1400
box -36 -19 303 1000
use PadBiDir  PadBiDir_10
timestamp 1711830429
transform 0 -1 -1500 -1 0 100
box -36 -19 303 1000
use PadBiDir  PadBiDir_11
timestamp 1711830429
transform 0 -1 -1500 1 0 400
box -36 -19 303 1000
use PadBiDir  PadBiDir_12
timestamp 1711830429
transform 0 -1 -1500 1 0 700
box -36 -19 303 1000
use PadBiDir  PadBiDir_13
timestamp 1711830429
transform 0 -1 -1500 1 0 1000
box -36 -19 303 1000
use PadBiDir  PadBiDir_14
timestamp 1711830429
transform 0 -1 -1500 1 0 1300
box -36 -19 303 1000
use PadBiDir  PadBiDir_15
timestamp 1711830429
transform 0 1 3300 1 0 100
box -36 -19 303 1000
use PadBiDir  PadBiDir_16
timestamp 1711830429
transform 0 1 3300 1 0 400
box -36 -19 303 1000
use PadBiDir  PadBiDir_17
timestamp 1711830429
transform 0 1 3300 1 0 700
box -36 -19 303 1000
use PadBiDir  PadBiDir_18
timestamp 1711830429
transform 0 1 3300 1 0 1000
box -36 -19 303 1000
use PadBiDir  PadBiDir_19
timestamp 1711830429
transform 0 1 3300 1 0 1300
box -36 -19 303 1000
use PadGnd  PadGnd_0
timestamp 1711831454
transform 0 -1 -1500 -1 0 400
box -3 -11 303 1000
use PadGnd  PadGnd_1
timestamp 1711831454
transform 0 1 3300 -1 0 100
box -3 -11 303 1000
use PadVdd  PadVdd_0
timestamp 1711831643
transform 1 0 2400 0 1 3400
box -3 -16 303 1000
use PadVdd  PadVdd_1
timestamp 1711831643
transform 1 0 1500 0 -1 -1400
box -3 -16 303 1000
use top_module  top_module_0
timestamp 1714281807
transform 1 0 -599 0 1 -492
box 0 0 3080 3040
<< end >>
