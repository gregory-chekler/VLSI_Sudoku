magic
tech scmos
timestamp 1711831643
<< nwell >>
rect 20 740 280 1000
rect 17 429 283 653
rect -3 248 303 330
rect -3 10 11 248
rect 289 10 303 248
rect -3 -4 303 10
<< pwell >>
rect -3 656 303 673
rect -3 426 14 656
rect 286 426 303 656
rect -3 340 303 426
rect 11 10 289 248
<< ntransistor >>
rect 38 215 138 218
rect 162 215 262 218
rect 38 170 138 173
rect 38 149 138 152
rect 162 170 262 173
rect 162 149 262 152
rect 38 105 138 108
rect 38 84 138 87
rect 162 105 262 108
rect 162 84 262 87
rect 38 40 138 43
rect 162 40 262 43
<< ndiffusion >>
rect 38 226 138 227
rect 38 222 41 226
rect 95 222 138 226
rect 38 218 138 222
rect 162 226 262 227
rect 162 222 205 226
rect 259 222 262 226
rect 162 218 262 222
rect 38 199 138 215
rect 38 195 56 199
rect 120 195 138 199
rect 38 193 138 195
rect 38 189 56 193
rect 120 189 138 193
rect 38 173 138 189
rect 38 166 138 170
rect 38 162 41 166
rect 120 162 138 166
rect 38 160 138 162
rect 38 156 41 160
rect 120 156 138 160
rect 38 152 138 156
rect 38 133 138 149
rect 38 124 56 133
rect 120 124 138 133
rect 38 108 138 124
rect 162 199 262 215
rect 162 195 180 199
rect 244 195 262 199
rect 162 193 262 195
rect 162 189 180 193
rect 244 189 262 193
rect 162 173 262 189
rect 162 166 262 170
rect 162 162 180 166
rect 259 162 262 166
rect 162 160 262 162
rect 162 156 180 160
rect 259 156 262 160
rect 162 152 262 156
rect 38 101 138 105
rect 38 97 41 101
rect 120 97 138 101
rect 38 95 138 97
rect 38 91 41 95
rect 120 91 138 95
rect 38 87 138 91
rect 38 68 138 84
rect 38 59 56 68
rect 120 59 138 68
rect 38 43 138 59
rect 162 133 262 149
rect 162 124 180 133
rect 244 124 262 133
rect 162 108 262 124
rect 162 101 262 105
rect 162 97 180 101
rect 259 97 262 101
rect 162 95 262 97
rect 162 91 180 95
rect 259 91 262 95
rect 162 87 262 91
rect 162 68 262 84
rect 162 59 180 68
rect 244 59 262 68
rect 162 43 262 59
rect 38 36 138 40
rect 38 32 41 36
rect 95 32 138 36
rect 38 31 138 32
rect 162 36 262 40
rect 162 32 205 36
rect 259 32 262 36
rect 162 31 262 32
<< ndcontact >>
rect 41 222 95 226
rect 205 222 259 226
rect 56 195 120 199
rect 56 189 120 193
rect 41 162 120 166
rect 41 156 120 160
rect 56 124 120 133
rect 180 195 244 199
rect 180 189 244 193
rect 180 162 259 166
rect 180 156 259 160
rect 41 97 120 101
rect 41 91 120 95
rect 56 59 120 68
rect 180 124 244 133
rect 180 97 259 101
rect 180 91 259 95
rect 180 59 244 68
rect 41 32 95 36
rect 205 32 259 36
<< psubstratepdiff >>
rect 0 669 300 670
rect 0 660 1 669
rect 95 660 204 669
rect 298 660 300 669
rect 0 659 300 660
rect 0 658 11 659
rect 0 424 1 658
rect 10 424 11 658
rect 289 658 300 659
rect 0 423 11 424
rect 289 424 290 658
rect 299 424 300 658
rect 289 423 300 424
rect 0 418 300 423
rect 0 414 143 418
rect 157 414 204 418
rect 298 414 300 418
rect 0 413 300 414
rect 0 409 2 413
rect 96 409 300 413
rect 0 408 300 409
rect 0 404 143 408
rect 157 404 204 408
rect 298 404 300 408
rect 0 403 300 404
rect 0 399 2 403
rect 96 399 300 403
rect 0 398 300 399
rect 0 394 143 398
rect 157 394 204 398
rect 298 394 300 398
rect 0 393 300 394
rect 0 389 2 393
rect 96 389 300 393
rect 0 388 300 389
rect 0 384 143 388
rect 157 384 204 388
rect 298 384 300 388
rect 0 383 300 384
rect 0 379 2 383
rect 96 379 300 383
rect 0 378 300 379
rect 0 374 143 378
rect 157 374 204 378
rect 298 374 300 378
rect 0 373 300 374
rect 0 369 2 373
rect 96 369 300 373
rect 0 368 300 369
rect 0 364 143 368
rect 157 364 204 368
rect 298 364 300 368
rect 0 363 300 364
rect 0 359 2 363
rect 96 359 300 363
rect 0 358 300 359
rect 0 354 143 358
rect 157 354 204 358
rect 298 354 300 358
rect 0 348 300 354
rect 0 344 2 348
rect 96 344 143 348
rect 157 344 204 348
rect 298 344 300 348
rect 0 343 300 344
rect 14 243 286 245
rect 14 240 202 243
rect 14 236 19 240
rect 98 236 202 240
rect 14 234 202 236
rect 281 234 286 243
rect 14 232 286 234
rect 14 28 24 232
rect 28 229 39 232
rect 28 29 30 229
rect 38 228 39 229
rect 98 229 202 232
rect 98 228 138 229
rect 38 227 138 228
rect 142 222 158 229
rect 142 218 145 222
rect 154 218 158 222
rect 162 228 202 229
rect 261 229 277 232
rect 261 228 262 229
rect 162 227 262 228
rect 142 214 158 218
rect 142 210 145 214
rect 154 210 158 214
rect 142 206 158 210
rect 142 202 145 206
rect 154 202 158 206
rect 142 134 158 202
rect 142 130 145 134
rect 154 130 158 134
rect 142 126 158 130
rect 142 122 145 126
rect 154 122 158 126
rect 142 62 158 122
rect 142 58 145 62
rect 154 58 158 62
rect 142 54 158 58
rect 142 50 145 54
rect 154 50 158 54
rect 142 46 158 50
rect 142 42 145 46
rect 154 42 158 46
rect 38 29 138 31
rect 142 38 158 42
rect 142 34 145 38
rect 154 34 158 38
rect 142 29 158 34
rect 162 29 262 31
rect 270 29 277 229
rect 28 28 277 29
rect 281 28 286 232
rect 14 26 286 28
rect 14 22 19 26
rect 98 22 202 26
rect 281 22 286 26
rect 14 13 286 22
<< nsubstratendiff >>
rect 20 649 280 650
rect 20 645 23 649
rect 277 645 280 649
rect 20 639 280 645
rect 20 635 23 639
rect 277 635 280 639
rect 20 629 280 635
rect 20 625 23 629
rect 277 625 280 629
rect 20 619 280 625
rect 20 615 23 619
rect 277 615 280 619
rect 20 609 280 615
rect 20 605 23 609
rect 277 605 280 609
rect 20 599 280 605
rect 20 595 23 599
rect 277 595 280 599
rect 20 589 280 595
rect 20 585 23 589
rect 277 585 280 589
rect 20 579 280 585
rect 20 575 23 579
rect 277 575 280 579
rect 20 569 280 575
rect 20 565 23 569
rect 277 565 280 569
rect 20 559 280 565
rect 20 555 23 559
rect 277 555 280 559
rect 20 549 280 555
rect 20 545 23 549
rect 277 545 280 549
rect 20 539 280 545
rect 20 535 23 539
rect 277 535 280 539
rect 20 529 280 535
rect 20 525 23 529
rect 277 525 280 529
rect 20 519 280 525
rect 20 515 23 519
rect 277 515 280 519
rect 20 509 280 515
rect 20 505 23 509
rect 277 505 280 509
rect 20 499 280 505
rect 20 495 23 499
rect 277 495 280 499
rect 20 489 280 495
rect 20 485 23 489
rect 277 485 280 489
rect 20 479 280 485
rect 20 475 23 479
rect 277 475 280 479
rect 20 469 280 475
rect 20 465 23 469
rect 277 465 280 469
rect 20 459 280 465
rect 20 455 23 459
rect 277 455 280 459
rect 20 449 280 455
rect 20 445 23 449
rect 277 445 280 449
rect 20 439 280 445
rect 20 435 23 439
rect 277 435 280 439
rect 20 432 280 435
rect 0 326 300 327
rect 0 322 3 326
rect 297 322 300 326
rect 0 316 300 322
rect 0 312 3 316
rect 297 312 300 316
rect 0 306 300 312
rect 0 302 3 306
rect 297 302 300 306
rect 0 296 300 302
rect 0 292 3 296
rect 297 292 300 296
rect 0 286 300 292
rect 0 282 3 286
rect 297 282 300 286
rect 0 276 300 282
rect 0 272 3 276
rect 297 272 300 276
rect 0 266 300 272
rect 0 262 3 266
rect 297 262 300 266
rect 0 256 300 262
rect 0 2 2 256
rect 6 252 8 256
rect 292 252 294 256
rect 6 251 294 252
rect 6 7 8 251
rect 292 7 294 251
rect 6 6 294 7
rect 6 2 8 6
rect 92 2 203 6
rect 292 2 294 6
rect 298 2 300 256
rect 0 -1 300 2
<< psubstratepcontact >>
rect 1 660 95 669
rect 204 660 298 669
rect 1 424 10 658
rect 290 424 299 658
rect 143 414 157 418
rect 204 414 298 418
rect 2 409 96 413
rect 143 404 157 408
rect 204 404 298 408
rect 2 399 96 403
rect 143 394 157 398
rect 204 394 298 398
rect 2 389 96 393
rect 143 384 157 388
rect 204 384 298 388
rect 2 379 96 383
rect 143 374 157 378
rect 204 374 298 378
rect 2 369 96 373
rect 143 364 157 368
rect 204 364 298 368
rect 2 359 96 363
rect 143 354 157 358
rect 204 354 298 358
rect 2 344 96 348
rect 143 344 157 348
rect 204 344 298 348
rect 19 236 98 240
rect 202 234 281 243
rect 24 28 28 232
rect 39 228 98 232
rect 145 218 154 222
rect 202 228 261 232
rect 145 210 154 214
rect 145 202 154 206
rect 145 130 154 134
rect 145 122 154 126
rect 145 58 154 62
rect 145 50 154 54
rect 145 42 154 46
rect 145 34 154 38
rect 277 28 281 232
rect 19 22 98 26
rect 202 22 281 26
<< nsubstratencontact >>
rect 23 645 277 649
rect 23 635 277 639
rect 23 625 277 629
rect 23 615 277 619
rect 23 605 277 609
rect 23 595 277 599
rect 23 585 277 589
rect 23 575 277 579
rect 23 565 277 569
rect 23 555 277 559
rect 23 545 277 549
rect 23 535 277 539
rect 23 525 277 529
rect 23 515 277 519
rect 23 505 277 509
rect 23 495 277 499
rect 23 485 277 489
rect 23 475 277 479
rect 23 465 277 469
rect 23 455 277 459
rect 23 445 277 449
rect 23 435 277 439
rect 3 322 297 326
rect 3 312 297 316
rect 3 302 297 306
rect 3 292 297 296
rect 3 282 297 286
rect 3 272 297 276
rect 3 262 297 266
rect 2 2 6 256
rect 8 252 292 256
rect 8 2 92 6
rect 203 2 292 6
rect 294 2 298 256
<< polysilicon >>
rect 6 713 21 716
rect 24 713 39 716
rect 12 701 15 713
rect 24 710 27 713
rect 36 710 39 713
rect 24 707 39 710
rect 24 701 27 707
rect 36 701 39 707
rect 42 713 45 716
rect 42 710 51 713
rect 42 701 45 710
rect 48 707 51 710
rect 54 707 57 716
rect 48 704 57 707
rect 54 701 57 704
rect 60 713 63 716
rect 60 710 69 713
rect 60 701 63 710
rect 66 707 69 710
rect 72 707 75 716
rect 66 704 75 707
rect 72 701 75 704
rect 78 713 93 716
rect 96 713 111 716
rect 78 710 81 713
rect 96 710 99 713
rect 108 710 111 713
rect 78 707 93 710
rect 96 707 111 710
rect 190 707 205 710
rect 78 704 81 707
rect 78 701 93 704
rect 96 701 99 707
rect 105 701 108 707
rect 190 695 193 707
rect 196 701 199 707
rect 202 695 205 707
rect 208 707 223 710
rect 208 698 211 707
rect 220 698 223 707
rect 226 707 241 710
rect 244 707 259 710
rect 262 707 277 710
rect 226 704 229 707
rect 226 701 241 704
rect 238 698 241 701
rect 250 698 253 707
rect 262 704 265 707
rect 262 701 277 704
rect 274 698 277 701
rect 208 695 223 698
rect 226 695 241 698
rect 244 695 259 698
rect 262 695 277 698
rect 51 688 66 691
rect 69 688 84 691
rect 87 688 102 691
rect 51 679 54 688
rect 69 685 72 688
rect 87 685 90 688
rect 69 682 84 685
rect 87 682 102 685
rect 69 679 72 682
rect 99 679 102 682
rect 51 676 66 679
rect 69 676 84 679
rect 87 676 102 679
rect 31 216 38 218
rect 31 42 32 216
rect 36 215 38 216
rect 138 215 140 218
rect 36 173 37 215
rect 160 215 162 218
rect 262 216 269 218
rect 262 215 264 216
rect 36 170 38 173
rect 138 170 140 173
rect 36 152 37 170
rect 36 149 38 152
rect 138 149 140 152
rect 36 108 37 149
rect 263 173 264 215
rect 160 170 162 173
rect 262 170 264 173
rect 263 152 264 170
rect 160 149 162 152
rect 262 149 264 152
rect 36 105 38 108
rect 138 105 140 108
rect 36 87 37 105
rect 36 84 38 87
rect 138 84 140 87
rect 36 43 37 84
rect 263 108 264 149
rect 160 105 162 108
rect 262 105 264 108
rect 263 87 264 105
rect 160 84 162 87
rect 262 84 264 87
rect 36 42 38 43
rect 31 40 38 42
rect 138 40 140 43
rect 263 43 264 84
rect 160 40 162 43
rect 262 42 264 43
rect 268 42 269 216
rect 262 40 269 42
<< polycontact >>
rect 32 42 36 216
rect 264 42 268 216
<< metal1 >>
rect 20 997 280 1000
rect 20 743 23 997
rect 277 743 280 997
rect 20 740 280 743
rect 62 730 238 740
rect 72 720 228 730
rect 82 710 218 720
rect 92 700 208 710
rect 0 669 99 670
rect 0 660 1 669
rect 95 660 99 669
rect 0 659 99 660
rect 0 658 10 659
rect 0 424 1 658
rect 102 650 198 700
rect 201 669 300 670
rect 201 660 204 669
rect 298 660 300 669
rect 201 659 300 660
rect 289 658 300 659
rect 50 649 280 650
rect 21 645 23 649
rect 277 645 280 649
rect 21 644 280 645
rect 21 640 23 644
rect 277 640 280 644
rect 21 639 280 640
rect 21 635 23 639
rect 277 635 280 639
rect 21 634 280 635
rect 21 630 23 634
rect 277 630 280 634
rect 21 629 280 630
rect 21 625 23 629
rect 277 625 280 629
rect 21 624 280 625
rect 21 620 23 624
rect 277 620 280 624
rect 21 619 280 620
rect 21 615 23 619
rect 277 615 280 619
rect 21 614 280 615
rect 21 610 23 614
rect 277 610 280 614
rect 21 609 280 610
rect 21 605 23 609
rect 277 605 280 609
rect 21 604 280 605
rect 21 600 23 604
rect 277 600 280 604
rect 21 599 280 600
rect 21 595 23 599
rect 277 595 280 599
rect 21 594 280 595
rect 21 590 23 594
rect 277 590 280 594
rect 21 589 280 590
rect 21 585 23 589
rect 277 585 280 589
rect 21 584 280 585
rect 21 580 23 584
rect 277 580 280 584
rect 21 579 280 580
rect 21 575 23 579
rect 277 575 280 579
rect 21 574 280 575
rect 21 570 23 574
rect 277 570 280 574
rect 21 569 280 570
rect 21 565 23 569
rect 277 565 280 569
rect 21 564 280 565
rect 21 560 23 564
rect 277 560 280 564
rect 21 559 280 560
rect 21 555 23 559
rect 277 555 280 559
rect 21 554 280 555
rect 21 550 23 554
rect 277 550 280 554
rect 21 549 280 550
rect 21 545 23 549
rect 277 545 280 549
rect 21 544 280 545
rect 21 540 23 544
rect 277 540 280 544
rect 21 539 280 540
rect 21 535 23 539
rect 277 535 280 539
rect 21 534 280 535
rect 21 530 23 534
rect 277 530 280 534
rect 21 529 280 530
rect 21 525 23 529
rect 277 525 280 529
rect 21 524 280 525
rect 21 520 23 524
rect 277 520 280 524
rect 21 519 280 520
rect 21 515 23 519
rect 277 515 280 519
rect 21 514 280 515
rect 21 510 23 514
rect 277 510 280 514
rect 21 509 280 510
rect 21 505 23 509
rect 277 505 280 509
rect 21 504 280 505
rect 21 500 23 504
rect 277 500 280 504
rect 21 499 280 500
rect 21 495 23 499
rect 277 495 280 499
rect 21 494 280 495
rect 21 490 23 494
rect 277 490 280 494
rect 21 489 280 490
rect 21 485 23 489
rect 277 485 280 489
rect 21 484 280 485
rect 21 480 23 484
rect 277 480 280 484
rect 21 479 280 480
rect 21 475 23 479
rect 277 475 280 479
rect 21 474 280 475
rect 21 470 23 474
rect 277 470 280 474
rect 21 469 280 470
rect 21 465 23 469
rect 277 465 280 469
rect 21 464 280 465
rect 21 460 23 464
rect 277 460 280 464
rect 21 459 280 460
rect 21 455 23 459
rect 277 455 280 459
rect 21 454 280 455
rect 21 450 23 454
rect 277 450 280 454
rect 21 449 280 450
rect 21 445 23 449
rect 277 445 280 449
rect 21 444 280 445
rect 21 440 23 444
rect 277 440 280 444
rect 21 439 280 440
rect 21 435 23 439
rect 277 435 280 439
rect 21 433 280 435
rect 0 419 10 424
rect 102 424 198 433
rect 0 418 99 419
rect 0 414 2 418
rect 96 414 99 418
rect 0 413 99 414
rect 0 409 2 413
rect 96 409 99 413
rect 0 408 99 409
rect 0 404 2 408
rect 96 404 99 408
rect 0 403 99 404
rect 0 399 2 403
rect 96 399 99 403
rect 0 398 99 399
rect 0 394 2 398
rect 96 394 99 398
rect 0 393 99 394
rect 0 389 2 393
rect 96 389 99 393
rect 0 388 99 389
rect 0 384 2 388
rect 96 384 99 388
rect 0 383 99 384
rect 0 379 2 383
rect 96 379 99 383
rect 0 378 99 379
rect 0 374 2 378
rect 96 374 99 378
rect 0 373 99 374
rect 0 369 2 373
rect 96 369 99 373
rect 0 368 99 369
rect 0 364 2 368
rect 96 364 99 368
rect 0 363 99 364
rect 0 359 2 363
rect 96 359 99 363
rect 0 358 99 359
rect 0 349 2 358
rect 96 349 99 358
rect 0 348 99 349
rect 0 344 2 348
rect 96 344 99 348
rect 102 340 140 424
rect 143 418 157 421
rect 143 413 157 414
rect 143 408 157 409
rect 143 403 157 404
rect 143 398 157 399
rect 143 393 157 394
rect 143 388 157 389
rect 143 383 157 384
rect 143 378 157 379
rect 143 373 157 374
rect 143 368 157 369
rect 143 363 157 364
rect 143 358 157 359
rect 143 353 157 354
rect 143 348 157 349
rect 160 340 198 424
rect 289 424 290 658
rect 299 424 300 658
rect 289 419 300 424
rect 201 418 300 419
rect 201 414 204 418
rect 298 414 300 418
rect 201 413 300 414
rect 201 409 204 413
rect 298 409 300 413
rect 201 408 300 409
rect 201 404 204 408
rect 298 404 300 408
rect 201 403 300 404
rect 201 399 204 403
rect 298 399 300 403
rect 201 398 300 399
rect 201 394 204 398
rect 298 394 300 398
rect 201 393 300 394
rect 201 389 204 393
rect 298 389 300 393
rect 201 388 300 389
rect 201 384 204 388
rect 298 384 300 388
rect 201 383 300 384
rect 201 379 204 383
rect 298 379 300 383
rect 201 378 300 379
rect 201 374 204 378
rect 298 374 300 378
rect 201 373 300 374
rect 201 369 204 373
rect 298 369 300 373
rect 201 368 300 369
rect 201 364 204 368
rect 298 364 300 368
rect 201 363 300 364
rect 201 359 204 363
rect 298 359 300 363
rect 201 358 300 359
rect 201 354 204 358
rect 298 354 300 358
rect 201 353 300 354
rect 201 349 204 353
rect 298 349 300 353
rect 201 348 300 349
rect 201 344 204 348
rect 298 344 300 348
rect 102 326 198 340
rect 0 322 3 326
rect 297 322 300 326
rect 0 321 300 322
rect 0 317 3 321
rect 297 317 300 321
rect 0 316 300 317
rect 0 312 3 316
rect 297 312 300 316
rect 0 311 300 312
rect 0 307 3 311
rect 297 307 300 311
rect 0 306 300 307
rect 0 302 3 306
rect 297 302 300 306
rect 0 301 300 302
rect 0 297 3 301
rect 297 297 300 301
rect 0 296 300 297
rect 0 292 3 296
rect 297 292 300 296
rect 0 291 300 292
rect 0 287 3 291
rect 297 287 300 291
rect 0 286 300 287
rect 0 282 3 286
rect 297 282 300 286
rect 0 281 300 282
rect 0 277 3 281
rect 297 277 300 281
rect 0 276 300 277
rect 0 272 3 276
rect 297 272 300 276
rect 0 271 300 272
rect 0 267 3 271
rect 297 267 300 271
rect 0 266 300 267
rect 0 262 3 266
rect 297 262 300 266
rect 0 261 300 262
rect 0 257 8 261
rect 292 257 300 261
rect 0 256 300 257
rect 0 2 2 256
rect 6 252 8 256
rect 292 252 294 256
rect 6 251 294 252
rect 6 7 8 251
rect 14 240 99 245
rect 14 236 19 240
rect 98 236 99 240
rect 14 232 99 236
rect 14 227 24 232
rect 14 28 19 227
rect 23 28 24 227
rect 28 228 39 232
rect 98 228 99 232
rect 28 226 99 228
rect 28 222 41 226
rect 95 222 99 226
rect 28 216 99 222
rect 28 42 32 216
rect 36 214 99 216
rect 36 195 39 214
rect 53 210 57 214
rect 96 210 99 214
rect 102 229 198 251
rect 102 207 142 229
rect 36 193 53 195
rect 36 174 39 193
rect 56 199 142 207
rect 157 207 198 229
rect 201 243 286 245
rect 201 234 202 243
rect 281 234 286 243
rect 201 232 286 234
rect 201 228 202 232
rect 261 228 277 232
rect 201 227 277 228
rect 201 226 272 227
rect 201 222 205 226
rect 259 222 272 226
rect 201 216 272 222
rect 201 214 264 216
rect 201 210 204 214
rect 243 210 247 214
rect 157 199 244 207
rect 120 195 180 199
rect 56 193 244 195
rect 120 189 180 193
rect 56 181 244 189
rect 261 195 264 214
rect 247 193 264 195
rect 53 174 57 178
rect 116 174 120 178
rect 36 166 120 174
rect 36 162 41 166
rect 36 160 120 162
rect 36 156 41 160
rect 36 148 120 156
rect 36 109 39 148
rect 53 144 57 148
rect 116 144 120 148
rect 123 141 177 181
rect 180 174 184 178
rect 243 174 247 178
rect 261 174 264 193
rect 180 166 264 174
rect 259 162 264 166
rect 180 160 264 162
rect 259 156 264 160
rect 180 148 264 156
rect 180 144 184 148
rect 243 144 247 148
rect 56 137 244 141
rect 56 133 142 137
rect 120 124 142 133
rect 56 119 142 124
rect 157 133 244 137
rect 157 124 180 133
rect 157 119 244 124
rect 56 116 244 119
rect 53 109 57 113
rect 116 109 120 113
rect 36 101 120 109
rect 36 97 41 101
rect 36 95 120 97
rect 36 91 41 95
rect 36 83 120 91
rect 36 44 39 83
rect 53 79 57 83
rect 116 79 120 83
rect 123 76 177 116
rect 180 109 184 113
rect 243 109 247 113
rect 261 109 264 148
rect 180 101 264 109
rect 259 97 264 101
rect 180 95 264 97
rect 259 91 264 95
rect 180 83 264 91
rect 180 79 184 83
rect 243 79 247 83
rect 56 69 244 76
rect 56 68 142 69
rect 120 59 142 68
rect 157 68 244 69
rect 56 51 142 59
rect 53 44 57 48
rect 96 44 99 48
rect 36 42 99 44
rect 28 36 99 42
rect 28 32 41 36
rect 95 32 99 36
rect 28 28 39 32
rect 98 28 99 32
rect 14 26 99 28
rect 14 22 19 26
rect 98 22 99 26
rect 14 21 99 22
rect 14 17 19 21
rect 98 17 99 21
rect 14 13 99 17
rect 102 27 142 51
rect 157 59 180 68
rect 157 51 244 59
rect 157 27 198 51
rect 6 6 99 7
rect 6 2 8 6
rect 92 2 99 6
rect 0 -1 99 2
rect 102 -1 198 27
rect 201 44 204 48
rect 243 44 247 48
rect 261 44 264 83
rect 201 42 264 44
rect 268 42 272 216
rect 201 36 272 42
rect 201 32 205 36
rect 259 32 272 36
rect 201 28 202 32
rect 261 28 272 32
rect 276 28 277 227
rect 281 28 286 232
rect 201 26 286 28
rect 201 22 202 26
rect 281 22 286 26
rect 201 21 286 22
rect 201 17 202 21
rect 281 17 286 21
rect 201 13 286 17
rect 292 7 294 251
rect 201 6 294 7
rect 201 2 203 6
rect 292 2 294 6
rect 298 2 300 256
rect 201 -1 300 2
rect 135 -16 158 -1
<< m2contact >>
rect 23 640 277 644
rect 23 630 277 634
rect 23 620 277 624
rect 23 610 277 614
rect 23 600 277 604
rect 23 590 277 594
rect 23 580 277 584
rect 23 570 277 574
rect 23 560 277 564
rect 23 550 277 554
rect 23 540 277 544
rect 23 530 277 534
rect 23 520 277 524
rect 23 510 277 514
rect 23 500 277 504
rect 23 490 277 494
rect 23 480 277 484
rect 23 470 277 474
rect 23 460 277 464
rect 23 450 277 454
rect 23 440 277 444
rect 2 414 96 418
rect 2 404 96 408
rect 2 394 96 398
rect 2 384 96 388
rect 2 374 96 378
rect 2 364 96 368
rect 2 349 96 358
rect 143 409 157 413
rect 143 399 157 403
rect 143 389 157 393
rect 143 379 157 383
rect 143 369 157 373
rect 143 359 157 363
rect 143 349 157 353
rect 204 409 298 413
rect 204 399 298 403
rect 204 389 298 393
rect 204 379 298 383
rect 204 369 298 373
rect 204 359 298 363
rect 204 349 298 353
rect 3 317 297 321
rect 3 307 297 311
rect 3 297 297 301
rect 3 287 297 291
rect 3 277 297 281
rect 3 267 297 271
rect 8 257 292 261
rect 19 28 23 227
rect 39 195 53 214
rect 57 210 96 214
rect 39 174 53 193
rect 145 222 154 226
rect 145 214 154 218
rect 145 206 154 210
rect 204 210 243 214
rect 247 195 261 214
rect 57 174 116 178
rect 39 109 53 148
rect 57 144 116 148
rect 184 174 243 178
rect 247 174 261 193
rect 184 144 243 148
rect 145 126 154 130
rect 57 109 116 113
rect 39 44 53 83
rect 57 79 116 83
rect 184 109 243 113
rect 247 109 261 148
rect 184 79 243 83
rect 57 44 96 48
rect 39 28 98 32
rect 19 17 98 21
rect 145 62 154 66
rect 145 54 154 58
rect 145 46 154 50
rect 145 38 154 42
rect 145 30 154 34
rect 204 44 243 48
rect 247 44 261 83
rect 202 28 261 32
rect 272 28 276 227
rect 202 17 281 21
<< metal2 >>
rect 20 997 280 1000
rect 20 743 23 997
rect 277 743 280 997
rect 20 740 280 743
rect 0 644 300 670
rect 0 640 23 644
rect 277 640 300 644
rect 0 634 300 640
rect 0 630 23 634
rect 277 630 300 634
rect 0 624 300 630
rect 0 620 23 624
rect 277 620 300 624
rect 0 614 300 620
rect 0 610 23 614
rect 277 610 300 614
rect 0 604 300 610
rect 0 600 23 604
rect 277 600 300 604
rect 0 594 300 600
rect 0 590 23 594
rect 277 590 300 594
rect 0 584 300 590
rect 0 580 23 584
rect 277 580 300 584
rect 0 574 300 580
rect 0 570 23 574
rect 277 570 300 574
rect 0 564 300 570
rect 0 560 23 564
rect 277 560 300 564
rect 0 554 300 560
rect 0 550 23 554
rect 277 550 300 554
rect 0 544 300 550
rect 0 540 23 544
rect 277 540 300 544
rect 0 534 300 540
rect 0 530 23 534
rect 277 530 300 534
rect 0 524 300 530
rect 0 520 23 524
rect 277 520 300 524
rect 0 514 300 520
rect 0 510 23 514
rect 277 510 300 514
rect 0 504 300 510
rect 0 500 23 504
rect 277 500 300 504
rect 0 494 300 500
rect 0 490 23 494
rect 277 490 300 494
rect 0 484 300 490
rect 0 480 23 484
rect 277 480 300 484
rect 0 474 300 480
rect 0 470 23 474
rect 277 470 300 474
rect 0 464 300 470
rect 0 460 23 464
rect 277 460 300 464
rect 0 454 300 460
rect 0 450 23 454
rect 277 450 300 454
rect 0 444 300 450
rect 0 440 23 444
rect 277 440 300 444
rect 0 418 300 424
rect 0 414 2 418
rect 96 414 300 418
rect 0 413 300 414
rect 0 409 143 413
rect 157 409 204 413
rect 298 409 300 413
rect 0 408 300 409
rect 0 404 2 408
rect 96 404 300 408
rect 0 403 300 404
rect 0 399 143 403
rect 157 399 204 403
rect 298 399 300 403
rect 0 398 300 399
rect 0 394 2 398
rect 96 394 300 398
rect 0 393 300 394
rect 0 389 143 393
rect 157 389 204 393
rect 298 389 300 393
rect 0 388 300 389
rect 0 384 2 388
rect 96 384 300 388
rect 0 383 300 384
rect 0 379 143 383
rect 157 379 204 383
rect 298 379 300 383
rect 0 378 300 379
rect 0 374 2 378
rect 96 374 300 378
rect 0 373 300 374
rect 0 369 143 373
rect 157 369 204 373
rect 298 369 300 373
rect 0 368 300 369
rect 0 364 2 368
rect 96 364 300 368
rect 0 363 300 364
rect 0 359 143 363
rect 157 359 204 363
rect 298 359 300 363
rect 0 358 300 359
rect 0 349 2 358
rect 96 353 300 358
rect 96 349 143 353
rect 157 349 204 353
rect 298 349 300 353
rect 0 344 300 349
rect 0 321 300 326
rect 0 317 3 321
rect 297 317 300 321
rect 0 311 300 317
rect 0 307 3 311
rect 297 307 300 311
rect 0 301 300 307
rect 0 297 3 301
rect 297 297 300 301
rect 0 291 300 297
rect 0 287 3 291
rect 297 287 300 291
rect 0 281 300 287
rect 0 277 3 281
rect 297 277 300 281
rect 0 271 300 277
rect 0 267 3 271
rect 297 267 300 271
rect 0 261 300 267
rect 0 257 8 261
rect 292 257 300 261
rect 0 246 300 257
rect 0 227 300 229
rect 0 28 19 227
rect 23 226 272 227
rect 23 222 145 226
rect 154 222 272 226
rect 23 218 272 222
rect 23 214 145 218
rect 154 214 272 218
rect 23 195 39 214
rect 53 210 57 214
rect 96 210 204 214
rect 243 210 247 214
rect 53 206 145 210
rect 154 206 247 210
rect 53 195 247 206
rect 261 195 272 214
rect 23 193 272 195
rect 23 174 39 193
rect 53 178 247 193
rect 53 174 57 178
rect 116 174 184 178
rect 243 174 247 178
rect 261 174 272 193
rect 23 148 272 174
rect 23 109 39 148
rect 53 144 57 148
rect 116 144 184 148
rect 243 144 247 148
rect 53 130 247 144
rect 53 126 145 130
rect 154 126 247 130
rect 53 113 247 126
rect 53 109 57 113
rect 116 109 184 113
rect 243 109 247 113
rect 261 109 272 148
rect 23 83 272 109
rect 23 44 39 83
rect 53 79 57 83
rect 116 79 184 83
rect 243 79 247 83
rect 53 66 247 79
rect 53 62 145 66
rect 154 62 247 66
rect 53 58 247 62
rect 53 54 145 58
rect 154 54 247 58
rect 53 50 247 54
rect 53 48 145 50
rect 53 44 57 48
rect 96 46 145 48
rect 154 48 247 50
rect 154 46 204 48
rect 96 44 204 46
rect 243 44 247 48
rect 261 44 272 83
rect 23 42 272 44
rect 23 38 145 42
rect 154 38 272 42
rect 23 34 272 38
rect 23 32 145 34
rect 23 28 39 32
rect 98 30 145 32
rect 154 32 272 34
rect 154 30 202 32
rect 98 28 202 30
rect 261 28 272 32
rect 276 28 300 227
rect 0 21 300 28
rect 0 17 19 21
rect 98 17 202 21
rect 281 17 300 21
rect 0 6 300 17
rect 0 -1 98 6
rect 202 -1 300 6
<< pad >>
rect 23 743 277 997
<< labels >>
rlabel metal1 150 -1 150 -1 8 Vdd!
rlabel metal1 150 -9 150 -9 1 Vdd!
<< end >>
