magic
tech scmos
timestamp 1714281807
<< m2contact >>
rect -2 -2 2 2
<< end >>
