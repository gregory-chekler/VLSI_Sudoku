magic
tech scmos
timestamp 1714281807
<< metal1 >>
rect 14 3007 3066 3027
rect 38 2983 3042 3003
rect 38 2967 3042 2973
rect 524 2943 541 2946
rect 724 2943 741 2946
rect 1802 2943 1844 2946
rect 2074 2943 2092 2946
rect 2226 2943 2260 2946
rect 2402 2943 2420 2946
rect 242 2926 245 2935
rect 258 2933 268 2936
rect 474 2933 508 2936
rect 642 2933 652 2936
rect 682 2933 708 2936
rect 842 2933 868 2936
rect 1154 2926 1157 2935
rect 1482 2926 1485 2935
rect 1532 2933 1565 2936
rect 1770 2933 1796 2936
rect 1852 2933 1877 2936
rect 2100 2933 2125 2936
rect 2268 2933 2293 2936
rect 2428 2933 2445 2936
rect 156 2923 181 2926
rect 212 2923 245 2926
rect 252 2923 276 2926
rect 356 2923 381 2926
rect 580 2923 605 2926
rect 780 2923 805 2926
rect 1148 2923 1157 2926
rect 1308 2923 1333 2926
rect 1364 2923 1373 2926
rect 1412 2923 1437 2926
rect 1468 2923 1485 2926
rect 1492 2923 1525 2926
rect 1700 2923 1725 2926
rect 1756 2923 1765 2926
rect 2012 2923 2021 2926
rect 2164 2923 2173 2926
rect 2276 2923 2285 2926
rect 2604 2923 2613 2926
rect 2708 2923 2717 2926
rect 2764 2923 2773 2926
rect 2812 2923 2837 2926
rect 292 2913 317 2916
rect 468 2913 493 2916
rect 676 2913 693 2916
rect 14 2867 3066 2873
rect 836 2823 861 2826
rect 1388 2823 1397 2826
rect 1468 2823 1477 2826
rect 276 2813 301 2816
rect 452 2813 461 2816
rect 506 2813 556 2816
rect 562 2813 621 2816
rect 636 2813 645 2816
rect 716 2813 765 2816
rect 772 2813 820 2816
rect 892 2813 949 2816
rect 1186 2813 1212 2816
rect 1356 2813 1365 2816
rect 1426 2813 1452 2816
rect 1524 2813 1557 2816
rect 1732 2813 1757 2816
rect 1788 2813 1797 2816
rect 1844 2813 1869 2816
rect 1900 2813 1909 2816
rect 1956 2813 1981 2816
rect 2012 2813 2021 2816
rect 2068 2813 2077 2816
rect 2098 2813 2116 2816
rect 2218 2813 2244 2816
rect 2284 2813 2309 2816
rect 2346 2813 2372 2816
rect 2412 2813 2437 2816
rect 2516 2813 2533 2816
rect 2572 2813 2589 2816
rect 2596 2813 2621 2816
rect 2708 2813 2732 2816
rect 2788 2813 2797 2816
rect 298 2805 301 2813
rect 410 2803 420 2806
rect 434 2803 444 2806
rect 466 2803 548 2806
rect 578 2803 588 2806
rect 674 2803 684 2806
rect 732 2803 764 2806
rect 930 2803 948 2806
rect 1034 2803 1068 2806
rect 1106 2803 1148 2806
rect 1362 2805 1365 2813
rect 1388 2803 1405 2806
rect 1482 2803 1500 2806
rect 1572 2803 1597 2806
rect 1794 2805 1797 2813
rect 1906 2805 1909 2813
rect 2018 2805 2021 2813
rect 2050 2803 2060 2806
rect 2586 2805 2589 2813
rect 2610 2803 2628 2806
rect 2700 2803 2717 2806
rect 2858 2803 2884 2806
rect 2634 2793 2692 2796
rect 2850 2793 2876 2796
rect 38 2767 3042 2773
rect 1602 2743 1620 2746
rect 236 2733 245 2736
rect 354 2726 357 2735
rect 564 2733 581 2736
rect 1354 2727 1357 2735
rect 1412 2733 1429 2736
rect 1628 2733 1645 2736
rect 1858 2733 1876 2736
rect 1946 2733 1964 2736
rect 2084 2733 2093 2736
rect 2148 2733 2165 2736
rect 2268 2733 2277 2736
rect 2282 2733 2292 2736
rect 340 2723 357 2726
rect 364 2723 380 2726
rect 468 2723 493 2726
rect 524 2723 533 2726
rect 570 2723 596 2726
rect 602 2723 612 2726
rect 636 2723 653 2726
rect 772 2723 780 2726
rect 804 2723 813 2726
rect 986 2723 1004 2726
rect 1146 2723 1156 2726
rect 1292 2723 1317 2726
rect 1348 2724 1357 2727
rect 2394 2726 2397 2735
rect 2402 2733 2420 2736
rect 2538 2733 2572 2736
rect 2690 2733 2724 2736
rect 2748 2733 2797 2736
rect 2828 2733 2853 2736
rect 2538 2726 2541 2733
rect 1364 2723 1373 2726
rect 1378 2723 1388 2726
rect 1426 2723 1460 2726
rect 1492 2723 1509 2726
rect 1532 2723 1565 2726
rect 1740 2723 1749 2726
rect 1754 2723 1772 2726
rect 1828 2723 1877 2726
rect 1898 2723 1972 2726
rect 2058 2723 2068 2726
rect 2124 2723 2165 2726
rect 2250 2723 2300 2726
rect 2378 2723 2397 2726
rect 2506 2723 2516 2726
rect 2530 2723 2541 2726
rect 2596 2723 2637 2726
rect 2690 2723 2732 2726
rect 2770 2723 2812 2726
rect 2826 2723 2877 2726
rect 1562 2716 1565 2723
rect 1562 2713 1572 2716
rect 1596 2713 1613 2716
rect 2084 2713 2093 2716
rect 2162 2706 2165 2723
rect 2748 2713 2757 2716
rect 1562 2703 1588 2706
rect 2162 2703 2196 2706
rect 14 2667 3066 2673
rect 2026 2633 2037 2636
rect 2634 2633 2644 2636
rect 226 2616 229 2626
rect 1324 2623 1357 2626
rect 132 2613 157 2616
rect 188 2613 197 2616
rect 204 2613 260 2616
rect 356 2613 381 2616
rect 476 2613 517 2616
rect 684 2613 693 2616
rect 722 2613 748 2616
rect 890 2613 900 2616
rect 972 2613 997 2616
rect 1028 2613 1061 2616
rect 1068 2613 1084 2616
rect 1188 2613 1197 2616
rect 1250 2613 1308 2616
rect 1380 2613 1412 2616
rect 1444 2613 1453 2616
rect 1668 2613 1716 2616
rect 1754 2613 1796 2616
rect 1884 2613 1909 2616
rect 1996 2613 2021 2616
rect 2034 2615 2037 2633
rect 2052 2623 2093 2626
rect 2196 2613 2205 2616
rect 2244 2613 2284 2616
rect 2322 2613 2372 2616
rect 2452 2613 2501 2616
rect 2666 2613 2700 2616
rect 2738 2613 2788 2616
rect 194 2605 197 2613
rect 210 2603 252 2606
rect 284 2603 317 2606
rect 490 2603 540 2606
rect 690 2605 693 2613
rect 754 2603 764 2606
rect 826 2603 852 2606
rect 1058 2605 1061 2613
rect 1180 2603 1189 2606
rect 1236 2603 1293 2606
rect 1570 2603 1580 2606
rect 1634 2603 1644 2606
rect 1954 2603 1972 2606
rect 2058 2603 2108 2606
rect 2188 2603 2213 2606
rect 2274 2603 2292 2606
rect 2402 2603 2444 2606
rect 2538 2603 2572 2606
rect 2658 2603 2708 2606
rect 2812 2603 2829 2606
rect 2834 2603 2852 2606
rect 1114 2593 1172 2596
rect 1202 2593 1228 2596
rect 2138 2593 2180 2596
rect 2410 2593 2436 2596
rect 38 2567 3042 2573
rect 938 2543 956 2546
rect 978 2543 1012 2546
rect 1034 2543 1068 2546
rect 1546 2543 1572 2546
rect 258 2533 276 2536
rect 474 2526 477 2535
rect 490 2533 508 2536
rect 546 2533 596 2536
rect 786 2527 789 2535
rect 914 2527 917 2535
rect 964 2533 1013 2536
rect 1020 2533 1037 2536
rect 1076 2533 1101 2536
rect 1490 2533 1508 2536
rect 1580 2533 1613 2536
rect 1722 2533 1732 2536
rect 188 2523 213 2526
rect 244 2523 277 2526
rect 314 2523 324 2526
rect 452 2523 477 2526
rect 484 2523 516 2526
rect 594 2523 604 2526
rect 724 2523 749 2526
rect 780 2524 789 2527
rect 852 2523 869 2526
rect 908 2524 917 2527
rect 1962 2526 1965 2535
rect 2266 2526 2269 2535
rect 2394 2526 2397 2535
rect 2530 2533 2540 2536
rect 2530 2526 2533 2533
rect 2794 2526 2797 2535
rect 2820 2533 2869 2536
rect 1140 2523 1149 2526
rect 1428 2523 1453 2526
rect 1490 2523 1516 2526
rect 1522 2523 1573 2526
rect 1730 2523 1740 2526
rect 1780 2523 1805 2526
rect 1884 2523 1909 2526
rect 1940 2523 1965 2526
rect 2012 2523 2021 2526
rect 2108 2523 2133 2526
rect 2204 2523 2229 2526
rect 2260 2523 2269 2526
rect 2276 2523 2285 2526
rect 2332 2523 2349 2526
rect 2388 2523 2397 2526
rect 2404 2523 2413 2526
rect 2468 2523 2485 2526
rect 2524 2523 2533 2526
rect 2538 2523 2548 2526
rect 2604 2523 2629 2526
rect 2700 2523 2725 2526
rect 2756 2523 2797 2526
rect 14 2467 3066 2473
rect 1524 2423 1557 2426
rect 2228 2423 2261 2426
rect 2356 2423 2365 2426
rect 2492 2423 2501 2426
rect 1554 2416 1557 2423
rect 338 2406 341 2416
rect 418 2413 436 2416
rect 588 2413 613 2416
rect 644 2413 669 2416
rect 1156 2413 1165 2416
rect 1268 2413 1277 2416
rect 1380 2413 1413 2416
rect 1442 2413 1508 2416
rect 1554 2413 1565 2416
rect 1756 2413 1781 2416
rect 1868 2413 1893 2416
rect 1954 2413 1964 2416
rect 2108 2413 2117 2416
rect 2138 2413 2212 2416
rect 2290 2413 2340 2416
rect 2546 2413 2604 2416
rect 2618 2413 2660 2416
rect 2666 2413 2700 2416
rect 292 2403 341 2406
rect 364 2403 397 2406
rect 418 2403 428 2406
rect 508 2403 549 2406
rect 666 2405 669 2413
rect 788 2403 853 2406
rect 860 2403 917 2406
rect 924 2403 957 2406
rect 1444 2403 1453 2406
rect 1572 2403 1605 2406
rect 1748 2403 1773 2406
rect 1778 2405 1781 2413
rect 1804 2403 1813 2406
rect 1980 2403 1989 2406
rect 2018 2403 2028 2406
rect 2058 2403 2100 2406
rect 2114 2405 2117 2413
rect 2140 2403 2149 2406
rect 2228 2403 2237 2406
rect 2378 2403 2404 2406
rect 2498 2403 2532 2406
rect 2620 2403 2629 2406
rect 2716 2403 2725 2406
rect 2780 2403 2797 2406
rect 458 2393 500 2396
rect 682 2393 708 2396
rect 738 2393 780 2396
rect 794 2393 852 2396
rect 874 2393 916 2396
rect 1706 2393 1740 2396
rect 2378 2393 2381 2403
rect 2498 2393 2501 2403
rect 2514 2393 2524 2396
rect 2722 2393 2772 2396
rect 38 2367 3042 2373
rect 370 2343 389 2346
rect 290 2326 293 2335
rect 364 2333 381 2336
rect 386 2326 389 2343
rect 458 2326 461 2345
rect 946 2343 964 2346
rect 1594 2343 1628 2346
rect 2090 2343 2116 2346
rect 468 2333 501 2336
rect 922 2333 972 2336
rect 1082 2333 1100 2336
rect 1130 2333 1148 2336
rect 1258 2333 1268 2336
rect 1322 2333 1364 2336
rect 1378 2333 1388 2336
rect 1842 2333 1860 2336
rect 1874 2326 1877 2335
rect 1964 2333 1989 2336
rect 2156 2333 2229 2336
rect 2666 2333 2692 2336
rect 2730 2333 2740 2336
rect 212 2323 237 2326
rect 268 2323 293 2326
rect 300 2323 357 2326
rect 386 2323 461 2326
rect 476 2323 485 2326
rect 540 2323 549 2326
rect 988 2323 1037 2326
rect 1108 2323 1125 2326
rect 1250 2323 1276 2326
rect 1300 2323 1365 2326
rect 1372 2323 1389 2326
rect 1396 2323 1405 2326
rect 1468 2323 1493 2326
rect 1538 2323 1556 2326
rect 1570 2323 1629 2326
rect 1780 2323 1789 2326
rect 1868 2323 1877 2326
rect 2084 2323 2101 2326
rect 2268 2323 2277 2326
rect 2436 2323 2461 2326
rect 2556 2323 2565 2326
rect 2604 2323 2629 2326
rect 2660 2323 2677 2326
rect 2700 2323 2748 2326
rect 1052 2313 1061 2316
rect 1076 2313 1093 2316
rect 1308 2313 1365 2316
rect 14 2267 3066 2273
rect 1066 2233 1132 2236
rect 1170 2233 1197 2236
rect 1012 2223 1029 2226
rect 1060 2223 1116 2226
rect 1146 2223 1188 2226
rect 300 2213 325 2216
rect 362 2213 404 2216
rect 418 2213 437 2216
rect 444 2213 477 2216
rect 684 2213 693 2216
rect 724 2213 733 2216
rect 772 2213 797 2216
rect 834 2213 852 2216
rect 924 2213 933 2216
rect 1010 2213 1052 2216
rect 1194 2215 1197 2233
rect 1212 2223 1245 2226
rect 1754 2223 1812 2226
rect 1836 2223 1845 2226
rect 1300 2213 1333 2216
rect 1356 2213 1381 2216
rect 1532 2213 1565 2216
rect 1722 2213 1748 2216
rect 1900 2213 1917 2216
rect 1980 2213 2005 2216
rect 2010 2213 2069 2216
rect 2108 2213 2125 2216
rect 2444 2213 2461 2216
rect 2548 2213 2573 2216
rect 2604 2213 2637 2216
rect 2706 2213 2757 2216
rect 2786 2213 2845 2216
rect 2892 2213 2901 2216
rect 2948 2213 2957 2216
rect 434 2205 437 2213
rect 2002 2206 2005 2213
rect 706 2203 716 2206
rect 874 2203 900 2206
rect 938 2203 988 2206
rect 1018 2203 1044 2206
rect 1306 2203 1348 2206
rect 1482 2203 1508 2206
rect 1556 2203 1628 2206
rect 1650 2203 1708 2206
rect 1730 2203 1740 2206
rect 1850 2203 1868 2206
rect 1916 2203 1933 2206
rect 1938 2203 1948 2206
rect 2002 2203 2028 2206
rect 2234 2203 2300 2206
rect 2610 2203 2644 2206
rect 2754 2205 2757 2213
rect 2780 2203 2805 2206
rect 2626 2193 2636 2196
rect 38 2167 3042 2173
rect 2050 2143 2092 2146
rect 2410 2143 2420 2146
rect 410 2133 436 2136
rect 460 2133 469 2136
rect 482 2133 500 2136
rect 522 2133 564 2136
rect 666 2133 676 2136
rect 748 2133 757 2136
rect 852 2133 861 2136
rect 1146 2133 1164 2136
rect 1188 2133 1197 2136
rect 1202 2133 1212 2136
rect 1314 2133 1348 2136
rect 586 2126 604 2127
rect 1626 2126 1629 2135
rect 1652 2133 1660 2136
rect 1754 2133 1772 2136
rect 1786 2133 1836 2136
rect 1860 2133 1869 2136
rect 1906 2133 1940 2136
rect 1956 2133 1965 2136
rect 1970 2133 2020 2136
rect 2100 2133 2117 2136
rect 2684 2133 2709 2136
rect 2722 2133 2732 2136
rect 2748 2133 2757 2136
rect 2794 2133 2812 2136
rect 2842 2133 2884 2136
rect 1906 2126 1909 2133
rect 236 2123 253 2126
rect 348 2123 373 2126
rect 404 2123 437 2126
rect 498 2123 508 2126
rect 572 2124 604 2126
rect 572 2123 589 2124
rect 684 2123 709 2126
rect 746 2123 804 2126
rect 810 2123 836 2126
rect 898 2123 908 2126
rect 1084 2123 1109 2126
rect 1140 2123 1149 2126
rect 1154 2123 1172 2126
rect 1210 2123 1261 2126
rect 1266 2123 1276 2126
rect 1308 2123 1333 2126
rect 1356 2123 1373 2126
rect 1412 2123 1421 2126
rect 1572 2123 1629 2126
rect 1668 2123 1701 2126
rect 1780 2123 1844 2126
rect 1884 2123 1909 2126
rect 2108 2123 2117 2126
rect 2156 2123 2165 2126
rect 2218 2123 2244 2126
rect 2436 2123 2452 2126
rect 2572 2123 2589 2126
rect 2786 2123 2804 2126
rect 2858 2123 2892 2126
rect 498 2116 501 2123
rect 1210 2116 1213 2123
rect 460 2113 501 2116
rect 516 2113 541 2116
rect 596 2113 605 2116
rect 692 2113 701 2116
rect 924 2113 949 2116
rect 1188 2113 1213 2116
rect 1508 2113 1517 2116
rect 1532 2113 1557 2116
rect 2266 2113 2284 2116
rect 2604 2113 2613 2116
rect 946 2106 949 2113
rect 578 2103 612 2106
rect 946 2103 965 2106
rect 986 2103 1020 2106
rect 1490 2103 1524 2106
rect 14 2067 3066 2073
rect 1730 2043 1749 2046
rect 1746 2036 1749 2043
rect 442 2033 500 2036
rect 514 2033 556 2036
rect 618 2033 644 2036
rect 1746 2033 1797 2036
rect 250 2016 253 2026
rect 426 2023 484 2026
rect 514 2023 540 2026
rect 618 2023 628 2026
rect 922 2023 941 2026
rect 1156 2023 1181 2026
rect 1196 2023 1221 2026
rect 1484 2023 1501 2026
rect 618 2016 621 2023
rect 938 2016 941 2023
rect 1178 2016 1181 2023
rect 1706 2016 1709 2025
rect 1730 2023 1788 2026
rect 250 2013 316 2016
rect 394 2006 397 2016
rect 570 2013 621 2016
rect 724 2013 749 2016
rect 938 2013 948 2016
rect 962 2013 972 2016
rect 994 2013 1004 2016
rect 1052 2013 1077 2016
rect 1114 2013 1140 2016
rect 1178 2013 1229 2016
rect 1236 2013 1261 2016
rect 1266 2006 1269 2014
rect 1314 2013 1356 2016
rect 1418 2013 1428 2016
rect 1476 2013 1493 2016
rect 1532 2013 1565 2016
rect 1596 2013 1629 2016
rect 1636 2013 1669 2016
rect 1706 2013 1724 2016
rect 1794 2015 1797 2033
rect 1812 2023 1837 2026
rect 2156 2023 2165 2026
rect 370 2005 397 2006
rect 370 2003 396 2005
rect 578 2003 604 2006
rect 954 2003 964 2006
rect 978 2003 996 2006
rect 1156 2003 1165 2006
rect 1194 2003 1228 2006
rect 1250 2003 1269 2006
rect 1292 2003 1301 2006
rect 1306 2003 1364 2006
rect 1402 2003 1420 2006
rect 1434 2003 1468 2006
rect 1482 2003 1524 2006
rect 1642 2003 1692 2006
rect 1706 2003 1716 2006
rect 1818 2003 1836 2006
rect 1898 2005 1901 2016
rect 1914 2013 1940 2016
rect 2010 2013 2036 2016
rect 2114 2013 2133 2016
rect 2228 2013 2237 2016
rect 2290 2013 2324 2016
rect 2362 2013 2428 2016
rect 2508 2013 2533 2016
rect 2564 2013 2589 2016
rect 2604 2013 2629 2016
rect 2708 2013 2748 2016
rect 2786 2013 2852 2016
rect 2866 2013 2884 2016
rect 2010 2006 2013 2013
rect 1938 2003 1948 2006
rect 1964 2003 2013 2006
rect 2018 2003 2044 2006
rect 2130 2005 2133 2013
rect 2362 2006 2365 2013
rect 2156 2003 2189 2006
rect 2298 2003 2332 2006
rect 2348 2003 2381 2006
rect 2444 2003 2453 2006
rect 2570 2003 2596 2006
rect 2626 2005 2629 2013
rect 2786 2006 2789 2013
rect 2722 2003 2756 2006
rect 2772 2003 2789 2006
rect 2802 2003 2844 2006
rect 2570 1993 2588 1996
rect 38 1967 3042 1973
rect 1994 1943 2036 1946
rect 2810 1943 2828 1946
rect 186 1926 189 1936
rect 250 1933 260 1936
rect 594 1933 636 1936
rect 186 1923 212 1926
rect 226 1923 268 1926
rect 314 1923 340 1926
rect 412 1923 421 1926
rect 532 1923 557 1926
rect 658 1923 661 1935
rect 722 1933 748 1936
rect 874 1933 900 1936
rect 924 1933 972 1936
rect 986 1933 1044 1936
rect 1074 1933 1084 1936
rect 1130 1935 1140 1936
rect 1130 1933 1141 1935
rect 1178 1933 1196 1936
rect 1250 1933 1277 1936
rect 1346 1933 1372 1936
rect 1410 1933 1436 1936
rect 1588 1933 1605 1936
rect 1810 1933 1820 1936
rect 1868 1933 1877 1936
rect 1898 1933 1964 1936
rect 2218 1933 2244 1936
rect 2396 1933 2421 1936
rect 1138 1926 1141 1933
rect 668 1923 677 1926
rect 772 1923 797 1926
rect 882 1923 908 1926
rect 1052 1923 1085 1926
rect 1092 1923 1141 1926
rect 1204 1923 1229 1926
rect 1244 1923 1261 1926
rect 1274 1925 1277 1933
rect 1874 1926 1877 1933
rect 2218 1926 2221 1933
rect 2538 1926 2541 1935
rect 2554 1933 2564 1936
rect 2770 1933 2796 1936
rect 2836 1933 2869 1936
rect 1314 1923 1364 1926
rect 1444 1923 1453 1926
rect 1874 1923 1885 1926
rect 1892 1923 1917 1926
rect 1972 1923 2021 1926
rect 2052 1923 2100 1926
rect 2148 1923 2173 1926
rect 2204 1923 2221 1926
rect 2268 1923 2309 1926
rect 2332 1923 2365 1926
rect 2516 1923 2541 1926
rect 2572 1923 2589 1926
rect 2652 1923 2677 1926
rect 2762 1923 2829 1926
rect 882 1916 885 1923
rect 276 1913 333 1916
rect 844 1913 885 1916
rect 988 1913 1005 1916
rect 1164 1913 1189 1916
rect 14 1867 3066 1873
rect 516 1823 541 1826
rect 676 1823 693 1826
rect 1036 1823 1045 1826
rect 1228 1823 1253 1826
rect 1308 1823 1341 1826
rect 124 1813 149 1816
rect 186 1813 204 1816
rect 380 1813 413 1816
rect 490 1813 549 1816
rect 570 1813 628 1816
rect 642 1813 660 1816
rect 802 1813 860 1816
rect 1010 1813 1020 1816
rect 1124 1813 1149 1816
rect 1180 1813 1213 1816
rect 1234 1813 1292 1816
rect 268 1803 285 1806
rect 410 1805 413 1813
rect 444 1803 477 1806
rect 538 1803 548 1806
rect 572 1803 581 1806
rect 634 1803 652 1806
rect 698 1803 732 1806
rect 762 1803 780 1806
rect 810 1803 852 1806
rect 890 1803 940 1806
rect 954 1803 996 1806
rect 1210 1805 1213 1813
rect 1338 1806 1341 1823
rect 1356 1813 1373 1816
rect 1476 1813 1485 1816
rect 1548 1813 1573 1816
rect 1604 1813 1629 1816
rect 1756 1813 1804 1816
rect 1258 1803 1284 1806
rect 1308 1803 1333 1806
rect 1338 1803 1348 1806
rect 1626 1805 1629 1813
rect 1850 1806 1853 1816
rect 1868 1813 1909 1816
rect 1786 1803 1796 1806
rect 1850 1803 1860 1806
rect 1906 1805 1909 1813
rect 1930 1806 1933 1826
rect 2020 1813 2045 1816
rect 2076 1813 2093 1816
rect 2252 1813 2316 1816
rect 2516 1813 2541 1816
rect 2572 1813 2581 1816
rect 2620 1813 2645 1816
rect 2676 1813 2709 1816
rect 2730 1813 2813 1816
rect 2956 1813 3013 1816
rect 1930 1803 1948 1806
rect 2122 1803 2140 1806
rect 2164 1803 2173 1806
rect 2290 1803 2324 1806
rect 2346 1803 2412 1806
rect 2738 1803 2748 1806
rect 2820 1803 2861 1806
rect 1666 1793 1740 1796
rect 2786 1793 2812 1796
rect 2786 1783 2789 1793
rect 38 1767 3042 1773
rect 2786 1743 2820 1746
rect 498 1733 532 1736
rect 556 1733 565 1736
rect 570 1733 628 1736
rect 892 1733 901 1736
rect 930 1733 940 1736
rect 970 1733 988 1736
rect 1058 1733 1092 1736
rect 1138 1733 1172 1736
rect 1186 1733 1196 1736
rect 1210 1733 1252 1736
rect 1546 1733 1556 1736
rect 1668 1733 1693 1736
rect 1764 1733 1797 1736
rect 2114 1733 2140 1736
rect 2468 1733 2493 1736
rect 2762 1733 2772 1736
rect 2828 1733 2861 1736
rect 1690 1726 1693 1733
rect 300 1723 325 1726
rect 370 1723 404 1726
rect 426 1723 484 1726
rect 490 1723 540 1726
rect 740 1723 765 1726
rect 802 1723 812 1726
rect 922 1723 948 1726
rect 1012 1723 1021 1726
rect 1162 1723 1180 1726
rect 1204 1723 1213 1726
rect 1260 1723 1277 1726
rect 1514 1723 1564 1726
rect 1676 1723 1685 1726
rect 1690 1723 1748 1726
rect 1940 1723 1965 1726
rect 2052 1723 2077 1726
rect 2108 1723 2125 1726
rect 2130 1723 2148 1726
rect 2274 1723 2333 1726
rect 2372 1723 2397 1726
rect 2588 1723 2597 1726
rect 2636 1723 2661 1726
rect 2692 1723 2701 1726
rect 2714 1723 2732 1726
rect 2746 1723 2821 1726
rect 556 1713 621 1716
rect 668 1713 693 1716
rect 964 1713 989 1716
rect 1268 1713 1285 1716
rect 1580 1713 1637 1716
rect 2164 1713 2189 1716
rect 650 1703 660 1706
rect 14 1667 3066 1673
rect 634 1633 645 1636
rect 634 1626 637 1633
rect 276 1623 309 1626
rect 532 1623 541 1626
rect 604 1623 637 1626
rect 644 1623 653 1626
rect 668 1623 709 1626
rect 948 1623 957 1626
rect 2004 1623 2021 1626
rect 154 1613 204 1616
rect 218 1613 268 1616
rect 490 1613 516 1616
rect 738 1613 749 1616
rect 764 1613 797 1616
rect 810 1613 820 1616
rect 890 1613 932 1616
rect 154 1603 157 1613
rect 282 1603 340 1606
rect 364 1603 420 1606
rect 452 1603 501 1606
rect 554 1603 580 1606
rect 674 1603 716 1606
rect 738 1605 741 1613
rect 994 1606 997 1614
rect 1084 1613 1093 1616
rect 1146 1613 1188 1616
rect 1242 1613 1268 1616
rect 1380 1613 1389 1616
rect 1394 1613 1445 1616
rect 1484 1613 1509 1616
rect 1548 1613 1573 1616
rect 1700 1613 1732 1616
rect 1764 1613 1805 1616
rect 1828 1613 1861 1616
rect 1900 1613 1981 1616
rect 2068 1613 2093 1616
rect 2180 1613 2205 1616
rect 2236 1613 2269 1616
rect 2284 1613 2349 1616
rect 2620 1613 2637 1616
rect 2778 1613 2821 1616
rect 1090 1606 1093 1613
rect 1386 1606 1389 1613
rect 746 1603 756 1606
rect 962 1603 997 1606
rect 1020 1603 1037 1606
rect 1090 1603 1108 1606
rect 1162 1603 1196 1606
rect 1218 1603 1260 1606
rect 1386 1603 1404 1606
rect 1442 1605 1445 1613
rect 1458 1603 1476 1606
rect 1660 1603 1669 1606
rect 1786 1603 1804 1606
rect 1898 1603 1940 1606
rect 1978 1605 1981 1613
rect 2050 1603 2060 1606
rect 2100 1603 2141 1606
rect 2242 1603 2276 1606
rect 2346 1605 2349 1613
rect 2372 1603 2389 1606
rect 2516 1603 2525 1606
rect 2668 1603 2677 1606
rect 2778 1603 2804 1606
rect 2828 1603 2869 1606
rect 962 1583 965 1603
rect 1858 1593 1884 1596
rect 2250 1593 2268 1596
rect 2490 1593 2508 1596
rect 1858 1583 1861 1593
rect 38 1567 3042 1573
rect 2386 1543 2412 1546
rect 298 1533 340 1536
rect 386 1533 396 1536
rect 410 1533 468 1536
rect 546 1533 580 1536
rect 618 1533 668 1536
rect 682 1533 724 1536
rect 932 1533 940 1536
rect 1074 1533 1132 1536
rect 1154 1533 1228 1536
rect 1250 1533 1300 1536
rect 1314 1533 1364 1536
rect 1386 1533 1460 1536
rect 212 1523 221 1526
rect 250 1523 268 1526
rect 348 1523 357 1526
rect 410 1515 413 1533
rect 418 1523 476 1526
rect 578 1523 588 1526
rect 618 1523 676 1526
rect 682 1516 685 1533
rect 1562 1526 1565 1535
rect 1618 1533 1660 1536
rect 2378 1533 2420 1536
rect 2516 1533 2525 1536
rect 2636 1533 2645 1536
rect 2724 1533 2773 1536
rect 706 1523 732 1526
rect 820 1523 829 1526
rect 876 1523 916 1526
rect 948 1523 957 1526
rect 962 1523 1020 1526
rect 1074 1523 1124 1526
rect 1156 1523 1165 1526
rect 1170 1523 1220 1526
rect 1308 1523 1349 1526
rect 1468 1523 1533 1526
rect 1548 1523 1565 1526
rect 1684 1523 1717 1526
rect 1780 1523 1797 1526
rect 1836 1523 1853 1526
rect 1948 1523 1957 1526
rect 1996 1523 2021 1526
rect 2260 1523 2277 1526
rect 2316 1523 2341 1526
rect 2372 1523 2405 1526
rect 2514 1523 2556 1526
rect 2562 1523 2620 1526
rect 2634 1523 2717 1526
rect 2868 1523 3013 1526
rect 682 1515 693 1516
rect 684 1513 693 1515
rect 962 1503 965 1523
rect 1162 1516 1165 1523
rect 1162 1513 1213 1516
rect 1588 1513 1645 1516
rect 2636 1513 2661 1516
rect 14 1467 3066 1473
rect 268 1423 309 1426
rect 412 1423 445 1426
rect 700 1423 741 1426
rect 1436 1423 1485 1426
rect 442 1416 445 1423
rect 164 1413 189 1416
rect 220 1413 253 1416
rect 260 1413 317 1416
rect 442 1413 485 1416
rect 492 1413 509 1416
rect 580 1413 597 1416
rect 658 1413 676 1416
rect 850 1413 868 1416
rect 908 1413 933 1416
rect 1020 1413 1029 1416
rect 1044 1413 1085 1416
rect 250 1405 253 1413
rect 1090 1406 1093 1414
rect 1130 1413 1196 1416
rect 1212 1413 1269 1416
rect 1418 1413 1428 1416
rect 1492 1413 1509 1416
rect 1556 1413 1565 1416
rect 1700 1413 1709 1416
rect 1722 1413 1732 1416
rect 1812 1413 1828 1416
rect 2012 1413 2020 1416
rect 2084 1413 2117 1416
rect 2260 1413 2325 1416
rect 2356 1413 2381 1416
rect 2420 1413 2445 1416
rect 2636 1413 2645 1416
rect 2692 1413 2717 1416
rect 1130 1406 1133 1413
rect 2714 1406 2717 1413
rect 2786 1413 2844 1416
rect 2786 1406 2789 1413
rect 298 1403 316 1406
rect 386 1403 396 1406
rect 466 1403 484 1406
rect 772 1403 781 1406
rect 842 1403 860 1406
rect 890 1403 900 1406
rect 922 1403 940 1406
rect 986 1403 996 1406
rect 1082 1403 1093 1406
rect 1116 1403 1133 1406
rect 1218 1403 1284 1406
rect 1386 1403 1420 1406
rect 1434 1403 1484 1406
rect 1548 1403 1565 1406
rect 1794 1403 1804 1406
rect 1810 1403 1820 1406
rect 1970 1403 1996 1406
rect 2050 1403 2076 1406
rect 2124 1403 2165 1406
rect 2290 1403 2348 1406
rect 2714 1403 2748 1406
rect 2764 1403 2789 1406
rect 2860 1403 2885 1406
rect 794 1393 820 1396
rect 1754 1393 1796 1396
rect 1962 1393 1988 1396
rect 2106 1393 2116 1396
rect 38 1367 3042 1373
rect 1634 1343 1644 1346
rect 2458 1343 2476 1346
rect 330 1333 340 1336
rect 634 1333 668 1336
rect 762 1333 788 1336
rect 804 1333 861 1336
rect 938 1333 972 1336
rect 1050 1333 1068 1336
rect 1396 1333 1413 1336
rect 1442 1333 1476 1336
rect 1594 1333 1652 1336
rect 1724 1333 1772 1336
rect 1788 1333 1821 1336
rect 1826 1333 1836 1336
rect 1860 1333 1885 1336
rect 2172 1333 2189 1336
rect 2378 1333 2420 1336
rect 2466 1333 2484 1336
rect 2546 1333 2556 1336
rect 2572 1333 2589 1336
rect 2658 1333 2676 1336
rect 938 1326 941 1333
rect 1546 1326 1564 1327
rect 1818 1326 1821 1333
rect 2586 1326 2589 1333
rect 252 1323 269 1326
rect 396 1323 421 1326
rect 460 1323 485 1326
rect 572 1323 597 1326
rect 642 1323 676 1326
rect 738 1323 780 1326
rect 812 1323 861 1326
rect 924 1323 941 1326
rect 996 1323 1005 1326
rect 1012 1323 1069 1326
rect 1082 1323 1148 1326
rect 1266 1323 1276 1326
rect 1298 1323 1324 1326
rect 1370 1323 1380 1326
rect 1428 1323 1437 1326
rect 1498 1324 1564 1326
rect 1498 1323 1549 1324
rect 1660 1323 1677 1326
rect 1796 1323 1805 1326
rect 1818 1323 1844 1326
rect 1924 1323 1949 1326
rect 1994 1323 2012 1326
rect 2026 1323 2044 1326
rect 2236 1323 2261 1326
rect 2292 1323 2309 1326
rect 2338 1323 2349 1326
rect 2356 1323 2365 1326
rect 2370 1323 2428 1326
rect 2492 1323 2541 1326
rect 2586 1323 2636 1326
rect 2700 1323 2741 1326
rect 2882 1323 2932 1326
rect 1084 1313 1125 1316
rect 1556 1313 1565 1316
rect 1580 1313 1629 1316
rect 2338 1315 2341 1323
rect 1626 1303 1629 1313
rect 2738 1306 2741 1323
rect 2748 1313 2757 1316
rect 2738 1303 2764 1306
rect 14 1267 3066 1273
rect 244 1223 253 1226
rect 132 1213 157 1216
rect 188 1213 229 1216
rect 258 1213 276 1216
rect 348 1213 373 1216
rect 482 1213 516 1216
rect 546 1213 596 1216
rect 626 1213 684 1216
rect 828 1213 861 1216
rect 868 1213 877 1216
rect 226 1205 229 1213
rect 292 1203 301 1206
rect 418 1203 436 1206
rect 474 1203 508 1206
rect 540 1203 565 1206
rect 834 1203 860 1206
rect 874 1195 877 1213
rect 890 1196 893 1214
rect 964 1213 989 1216
rect 1010 1213 1044 1216
rect 1010 1206 1013 1213
rect 996 1203 1013 1206
rect 1090 1206 1093 1236
rect 1650 1233 1708 1236
rect 2458 1226 2461 1246
rect 1116 1223 1125 1226
rect 1682 1216 1685 1226
rect 1692 1223 1701 1226
rect 2012 1223 2053 1226
rect 2452 1223 2461 1226
rect 1108 1213 1117 1216
rect 1162 1213 1172 1216
rect 1258 1213 1284 1216
rect 1356 1213 1381 1216
rect 1442 1213 1452 1216
rect 1548 1213 1565 1216
rect 1644 1213 1685 1216
rect 1772 1213 1828 1216
rect 1940 1213 1989 1216
rect 2100 1213 2117 1216
rect 2156 1213 2189 1216
rect 2220 1213 2284 1216
rect 1090 1203 1100 1206
rect 1130 1203 1164 1206
rect 1434 1203 1444 1206
rect 1476 1203 1493 1206
rect 1610 1203 1636 1206
rect 1810 1203 1836 1206
rect 1858 1203 1932 1206
rect 1986 1205 1989 1213
rect 2314 1206 2317 1214
rect 2322 1213 2365 1216
rect 2388 1213 2436 1216
rect 2620 1213 2645 1216
rect 2676 1213 2685 1216
rect 2698 1213 2740 1216
rect 2778 1213 2836 1216
rect 2850 1213 2884 1216
rect 2012 1203 2021 1206
rect 2170 1203 2196 1206
rect 2314 1203 2325 1206
rect 2362 1205 2365 1213
rect 2516 1203 2525 1206
rect 2530 1203 2548 1206
rect 2682 1205 2685 1213
rect 2778 1206 2781 1213
rect 2764 1203 2781 1206
rect 2794 1203 2828 1206
rect 2852 1203 2861 1206
rect 890 1193 940 1196
rect 970 1193 988 1196
rect 1810 1193 1813 1203
rect 2322 1193 2325 1203
rect 2498 1193 2508 1196
rect 38 1167 3042 1173
rect 770 1143 796 1146
rect 922 1143 948 1146
rect 1258 1143 1292 1146
rect 1498 1143 1548 1146
rect 234 1133 276 1136
rect 474 1126 477 1135
rect 506 1133 532 1136
rect 602 1133 620 1136
rect 706 1133 740 1136
rect 506 1126 509 1133
rect 452 1123 477 1126
rect 484 1123 509 1126
rect 530 1123 540 1126
rect 594 1123 628 1126
rect 722 1123 748 1126
rect 770 1116 773 1143
rect 804 1133 845 1136
rect 922 1126 925 1143
rect 1562 1136 1565 1146
rect 1986 1143 1996 1146
rect 2858 1143 2884 1146
rect 938 1133 956 1136
rect 1036 1133 1068 1136
rect 1090 1133 1116 1136
rect 1178 1133 1188 1136
rect 1210 1133 1244 1136
rect 1300 1133 1317 1136
rect 1404 1133 1428 1136
rect 1556 1133 1565 1136
rect 1650 1133 1700 1136
rect 1716 1133 1757 1136
rect 1852 1133 1877 1136
rect 2004 1133 2021 1136
rect 2164 1133 2173 1136
rect 2178 1133 2204 1136
rect 2226 1133 2285 1136
rect 2308 1133 2325 1136
rect 2330 1133 2340 1136
rect 2364 1133 2373 1136
rect 2818 1133 2844 1136
rect 2882 1133 2892 1136
rect 818 1123 868 1126
rect 884 1123 925 1126
rect 978 1123 1012 1126
rect 1066 1123 1076 1126
rect 1124 1123 1141 1126
rect 1196 1123 1245 1126
rect 1252 1123 1261 1126
rect 1380 1123 1413 1126
rect 1436 1123 1445 1126
rect 1650 1123 1653 1133
rect 1724 1123 1741 1126
rect 1788 1123 1821 1126
rect 1916 1123 1941 1126
rect 2060 1123 2069 1126
rect 2116 1123 2133 1126
rect 2282 1125 2285 1133
rect 2322 1126 2325 1133
rect 2322 1123 2348 1126
rect 676 1113 685 1116
rect 756 1113 773 1116
rect 1458 1113 1468 1116
rect 1636 1113 1685 1116
rect 2164 1113 2189 1116
rect 2370 1103 2373 1133
rect 2404 1123 2413 1126
rect 2460 1123 2469 1126
rect 2620 1123 2645 1126
rect 2756 1123 2781 1126
rect 2812 1123 2829 1126
rect 2882 1123 2885 1133
rect 14 1067 3066 1073
rect 658 1023 677 1026
rect 1180 1023 1221 1026
rect 2764 1023 2773 1026
rect 276 1013 285 1016
rect 452 1013 469 1016
rect 476 1013 525 1016
rect 562 1013 612 1016
rect 658 1013 661 1023
rect 698 1013 708 1016
rect 956 1013 973 1016
rect 1060 1013 1085 1016
rect 466 1005 469 1013
rect 522 1005 525 1013
rect 1106 1006 1109 1014
rect 1114 1013 1164 1016
rect 1218 1013 1228 1016
rect 1364 1013 1373 1016
rect 1452 1013 1477 1016
rect 1514 1013 1540 1016
rect 1612 1013 1637 1016
rect 1668 1013 1677 1016
rect 1684 1013 1701 1016
rect 1788 1013 1828 1016
rect 1972 1013 1989 1016
rect 2034 1013 2060 1016
rect 2148 1013 2173 1016
rect 2204 1013 2221 1016
rect 2284 1013 2293 1016
rect 2340 1013 2381 1016
rect 2388 1013 2421 1016
rect 2564 1013 2573 1016
rect 2708 1013 2741 1016
rect 2860 1013 2885 1016
rect 2916 1013 3013 1016
rect 794 1003 876 1006
rect 1018 1003 1052 1006
rect 1106 1003 1156 1006
rect 1180 1003 1229 1006
rect 1252 1003 1269 1006
rect 1370 1005 1373 1013
rect 1674 1005 1677 1013
rect 2100 1003 2109 1006
rect 2218 1005 2221 1013
rect 2378 1005 2381 1013
rect 2428 1003 2469 1006
rect 2588 1003 2613 1006
rect 850 993 868 996
rect 1066 993 1092 996
rect 1266 983 1269 1003
rect 1754 993 1772 996
rect 38 967 3042 973
rect 554 943 604 946
rect 434 933 500 936
rect 612 933 645 936
rect 650 926 653 935
rect 674 933 708 936
rect 730 933 772 936
rect 812 933 853 936
rect 290 923 332 926
rect 290 913 293 923
rect 378 913 404 916
rect 410 906 413 925
rect 482 923 508 926
rect 530 923 548 926
rect 626 923 653 926
rect 866 925 869 946
rect 1666 943 1676 946
rect 1994 943 2036 946
rect 2786 943 2796 946
rect 1644 933 1653 936
rect 1962 926 1965 935
rect 2044 933 2077 936
rect 2218 933 2252 936
rect 2738 933 2764 936
rect 2804 933 2845 936
rect 2738 926 2741 933
rect 1036 923 1061 926
rect 1348 923 1373 926
rect 1404 923 1413 926
rect 1418 923 1452 926
rect 1474 923 1508 926
rect 1554 923 1564 926
rect 1620 923 1629 926
rect 1692 923 1701 926
rect 1764 923 1781 926
rect 1820 923 1837 926
rect 1842 923 1868 926
rect 1940 923 1965 926
rect 2172 923 2229 926
rect 2340 923 2365 926
rect 2396 923 2437 926
rect 2466 923 2484 926
rect 2676 923 2701 926
rect 2732 923 2741 926
rect 2746 923 2797 926
rect 530 916 533 923
rect 516 913 533 916
rect 834 913 860 916
rect 906 913 932 916
rect 956 913 965 916
rect 1468 913 1501 916
rect 1884 913 1893 916
rect 1988 913 2029 916
rect 394 903 413 906
rect 826 903 876 906
rect 890 903 948 906
rect 14 867 3066 873
rect 1298 833 1332 836
rect 1132 823 1173 826
rect 1298 823 1316 826
rect 1340 823 1373 826
rect 2316 823 2333 826
rect 1298 816 1301 823
rect 268 813 293 816
rect 380 813 397 816
rect 572 813 581 816
rect 668 813 693 816
rect 764 813 789 816
rect 860 813 877 816
rect 1004 813 1029 816
rect 1060 813 1069 816
rect 1076 813 1085 816
rect 1098 813 1116 816
rect 1170 813 1180 816
rect 1212 813 1229 816
rect 1268 813 1301 816
rect 1066 805 1069 813
rect 1082 806 1085 813
rect 1082 803 1108 806
rect 1178 803 1188 806
rect 1210 803 1244 806
rect 1370 796 1373 823
rect 1378 803 1388 806
rect 1394 803 1397 814
rect 1444 813 1477 816
rect 1612 813 1621 816
rect 1660 813 1685 816
rect 1836 813 1861 816
rect 1898 813 1957 816
rect 2100 813 2109 816
rect 2148 813 2173 816
rect 2204 813 2221 816
rect 2252 814 2261 816
rect 2250 813 2261 814
rect 2266 813 2300 816
rect 2628 813 2677 816
rect 2706 813 2756 816
rect 2250 806 2253 813
rect 1410 803 1436 806
rect 1484 803 1517 806
rect 1722 803 1756 806
rect 1898 803 1924 806
rect 1964 803 2005 806
rect 2226 803 2244 806
rect 2250 803 2292 806
rect 2492 803 2533 806
rect 2650 803 2676 806
rect 2772 803 2797 806
rect 2828 803 2853 806
rect 1370 793 1380 796
rect 1450 793 1476 796
rect 2466 793 2484 796
rect 2786 793 2820 796
rect 38 767 3042 773
rect 290 743 340 746
rect 386 743 404 746
rect 514 743 572 746
rect 642 743 684 746
rect 762 743 796 746
rect 1034 743 1044 746
rect 1666 743 1676 746
rect 1994 743 2036 746
rect 2282 743 2308 746
rect 2506 743 2524 746
rect 290 733 348 736
rect 386 726 389 743
rect 394 733 412 736
rect 450 733 460 736
rect 474 733 508 736
rect 714 733 740 736
rect 786 733 804 736
rect 810 733 852 736
rect 1010 733 1052 736
rect 1154 733 1180 736
rect 1196 733 1205 736
rect 1346 726 1349 735
rect 1378 726 1381 735
rect 1404 733 1413 736
rect 1444 733 1461 736
rect 1658 733 1684 736
rect 1698 733 1708 736
rect 1922 733 1948 736
rect 1962 727 1965 735
rect 2044 733 2069 736
rect 2316 733 2333 736
rect 2500 733 2509 736
rect 2532 733 2565 736
rect 2866 733 2876 736
rect 266 723 284 726
rect 364 723 389 726
rect 420 723 461 726
rect 516 723 565 726
rect 588 723 628 726
rect 700 723 709 726
rect 756 723 797 726
rect 948 723 973 726
rect 1060 723 1085 726
rect 1204 723 1221 726
rect 1276 723 1301 726
rect 1332 723 1349 726
rect 1356 723 1381 726
rect 1596 723 1613 726
rect 1692 723 1725 726
rect 1764 723 1781 726
rect 1860 723 1869 726
rect 1916 723 1933 726
rect 1956 724 1965 727
rect 2212 723 2229 726
rect 2268 723 2309 726
rect 2458 723 2484 726
rect 2858 723 2884 726
rect 266 715 269 723
rect 1116 713 1165 716
rect 1404 713 1421 716
rect 14 667 3066 673
rect 1178 633 1197 636
rect 580 623 637 626
rect 652 623 685 626
rect 682 616 685 623
rect 1178 616 1181 633
rect 268 613 277 616
rect 324 613 349 616
rect 388 613 413 616
rect 500 613 509 616
rect 562 613 572 616
rect 610 613 644 616
rect 682 613 741 616
rect 762 613 804 616
rect 996 613 1021 616
rect 1052 613 1085 616
rect 1092 613 1117 616
rect 1140 613 1181 616
rect 1194 615 1197 633
rect 1212 623 1237 626
rect 1428 623 1437 626
rect 2044 623 2053 626
rect 2428 623 2445 626
rect 1284 613 1309 616
rect 1340 613 1365 616
rect 1372 613 1405 616
rect 1770 613 1788 616
rect 1924 613 1949 616
rect 2252 613 2293 616
rect 2300 613 2317 616
rect 2338 613 2412 616
rect 2484 613 2509 616
rect 2546 613 2556 616
rect 2674 613 2725 616
rect 2868 613 2989 616
rect 492 603 501 606
rect 546 603 564 606
rect 650 603 692 606
rect 738 595 741 613
rect 748 603 789 606
rect 1082 605 1085 613
rect 1114 605 1117 613
rect 1362 605 1365 613
rect 1402 605 1405 613
rect 1428 603 1445 606
rect 1476 603 1509 606
rect 1644 603 1653 606
rect 1804 603 1845 606
rect 1852 603 1869 606
rect 2116 603 2157 606
rect 2258 603 2292 606
rect 2314 605 2317 613
rect 2732 603 2773 606
rect 1610 593 1636 596
rect 1810 593 1844 596
rect 2074 593 2108 596
rect 38 567 3042 573
rect 460 543 508 546
rect 866 543 892 546
rect 1466 543 1476 546
rect 2194 536 2197 546
rect 2602 536 2605 546
rect 394 533 444 536
rect 516 533 557 536
rect 658 533 700 536
rect 858 533 900 536
rect 1058 533 1084 536
rect 1098 533 1132 536
rect 1370 526 1373 535
rect 1402 526 1405 535
rect 1428 533 1437 536
rect 1484 533 1517 536
rect 1674 526 1677 535
rect 2026 533 2044 536
rect 2114 526 2117 534
rect 2122 533 2164 536
rect 2194 533 2212 536
rect 2498 526 2501 534
rect 2564 533 2605 536
rect 2708 533 2756 536
rect 2778 533 2836 536
rect 2860 533 2869 536
rect 332 523 357 526
rect 596 523 605 526
rect 652 523 701 526
rect 796 523 821 526
rect 852 523 877 526
rect 908 523 949 526
rect 1156 523 1189 526
rect 1228 523 1253 526
rect 1292 523 1317 526
rect 1348 523 1373 526
rect 1380 523 1405 526
rect 1612 523 1629 526
rect 1652 523 1677 526
rect 1836 523 1853 526
rect 1956 523 1981 526
rect 2018 523 2052 526
rect 2066 523 2100 526
rect 2114 523 2165 526
rect 2300 523 2325 526
rect 2412 523 2429 526
rect 2468 523 2501 526
rect 2636 523 2661 526
rect 2690 523 2748 526
rect 2826 523 2844 526
rect 2858 523 2884 526
rect 698 513 701 523
rect 1700 513 1757 516
rect 14 467 3066 473
rect 2698 433 2717 436
rect 660 423 685 426
rect 1076 423 1125 426
rect 2652 423 2661 426
rect 260 413 269 416
rect 316 413 333 416
rect 354 413 364 416
rect 370 413 404 416
rect 538 413 573 416
rect 596 413 645 416
rect 828 413 853 416
rect 884 413 893 416
rect 940 413 965 416
rect 378 403 396 406
rect 420 403 429 406
rect 500 403 509 406
rect 570 405 573 413
rect 642 405 645 413
rect 1026 405 1029 416
rect 1036 413 1045 416
rect 1164 413 1197 416
rect 1228 413 1268 416
rect 1300 413 1333 416
rect 1492 413 1532 416
rect 1620 413 1645 416
rect 1820 413 1837 416
rect 1956 413 1996 416
rect 2042 413 2084 416
rect 1042 406 1045 413
rect 2394 406 2397 414
rect 2402 413 2460 416
rect 2498 413 2532 416
rect 2564 413 2589 416
rect 2620 413 2660 416
rect 2698 406 2701 433
rect 2762 413 2804 416
rect 2900 413 2933 416
rect 1042 403 1052 406
rect 1076 403 1085 406
rect 1380 403 1420 406
rect 1442 403 1468 406
rect 1690 403 1700 406
rect 1780 403 1789 406
rect 1842 403 1884 406
rect 1900 403 1909 406
rect 1922 403 1932 406
rect 2020 403 2045 406
rect 2266 403 2276 406
rect 2292 403 2301 406
rect 2314 403 2348 406
rect 2394 403 2453 406
rect 2458 403 2468 406
rect 2556 403 2565 406
rect 2570 403 2596 406
rect 2698 403 2732 406
rect 2834 403 2876 406
rect 1730 393 1772 396
rect 1786 393 1789 403
rect 38 367 3042 373
rect 442 343 477 346
rect 1130 343 1141 346
rect 474 336 477 343
rect 1138 336 1141 343
rect 228 333 293 336
rect 322 333 380 336
rect 394 333 412 336
rect 426 333 469 336
rect 474 333 484 336
rect 516 333 549 336
rect 658 333 684 336
rect 810 333 828 336
rect 842 333 876 336
rect 1010 333 1044 336
rect 1074 333 1100 336
rect 1124 333 1133 336
rect 1138 333 1181 336
rect 1204 333 1213 336
rect 1218 333 1268 336
rect 1292 333 1301 336
rect 1314 333 1324 336
rect 1378 333 1412 336
rect 1436 333 1453 336
rect 236 323 285 326
rect 290 325 293 333
rect 394 326 397 333
rect 466 326 469 333
rect 324 323 349 326
rect 388 323 397 326
rect 428 323 461 326
rect 466 323 492 326
rect 786 323 836 326
rect 866 323 884 326
rect 948 323 973 326
rect 1004 323 1021 326
rect 1052 323 1061 326
rect 1066 323 1108 326
rect 1178 325 1181 333
rect 1522 326 1525 335
rect 1674 333 1684 336
rect 1842 333 1860 336
rect 1884 333 1893 336
rect 2020 333 2037 336
rect 1610 326 1628 327
rect 1842 326 1845 333
rect 2042 326 2045 335
rect 2082 333 2100 336
rect 2124 333 2149 336
rect 2154 326 2157 335
rect 2274 333 2292 336
rect 2316 333 2325 336
rect 2402 333 2412 336
rect 2466 333 2492 336
rect 2516 333 2525 336
rect 2596 333 2605 336
rect 2692 333 2701 336
rect 2706 333 2740 336
rect 2764 333 2773 336
rect 2852 333 2869 336
rect 2466 326 2469 333
rect 1212 323 1269 326
rect 1348 323 1413 326
rect 1434 323 1508 326
rect 1522 323 1541 326
rect 1564 323 1573 326
rect 1594 324 1628 326
rect 1594 323 1613 324
rect 1658 323 1692 326
rect 1756 323 1789 326
rect 1818 323 1845 326
rect 2034 323 2045 326
rect 2130 323 2157 326
rect 2180 323 2189 326
rect 2244 323 2269 326
rect 2442 323 2469 326
rect 2490 323 2500 326
rect 2514 323 2580 326
rect 2762 323 2836 326
rect 2850 323 2884 326
rect 866 316 869 323
rect 538 313 556 316
rect 652 313 677 316
rect 844 313 869 316
rect 1124 313 1173 316
rect 1436 313 1445 316
rect 1594 313 1620 316
rect 1644 313 1669 316
rect 1708 313 1725 316
rect 546 303 572 306
rect 618 303 644 306
rect 1610 303 1636 306
rect 2034 293 2037 323
rect 2068 313 2093 316
rect 2372 313 2381 316
rect 14 267 3066 273
rect 922 253 957 256
rect 354 233 380 236
rect 300 213 325 216
rect 354 206 357 233
rect 388 223 413 226
rect 588 223 637 226
rect 292 203 357 206
rect 410 206 413 223
rect 866 216 869 226
rect 2402 216 2405 236
rect 418 213 436 216
rect 514 213 580 216
rect 586 213 677 216
rect 772 213 869 216
rect 1012 213 1045 216
rect 1092 213 1109 216
rect 1148 213 1173 216
rect 1276 213 1301 216
rect 1412 213 1437 216
rect 1468 213 1477 216
rect 1498 213 1516 216
rect 1676 213 1701 216
rect 1732 213 1757 216
rect 1876 213 1893 216
rect 1988 213 2013 216
rect 2044 213 2069 216
rect 2076 213 2085 216
rect 2226 213 2252 216
rect 2292 213 2317 216
rect 2348 213 2357 216
rect 2402 213 2429 216
rect 2468 213 2493 216
rect 2564 213 2589 216
rect 2620 213 2629 216
rect 2650 213 2709 216
rect 2748 213 2773 216
rect 410 203 428 206
rect 516 203 525 206
rect 586 203 644 206
rect 658 203 676 206
rect 690 203 756 206
rect 978 203 1004 206
rect 1170 205 1173 213
rect 1754 205 1757 213
rect 2066 205 2069 213
rect 2234 203 2244 206
rect 2402 203 2412 206
rect 2626 205 2629 213
rect 2860 203 2901 206
rect 258 193 284 196
rect 658 183 661 203
rect 772 193 781 196
rect 978 193 981 203
rect 38 167 3042 173
rect 828 143 837 146
rect 1346 143 1364 146
rect 1514 143 1532 146
rect 1674 143 1692 146
rect 1842 143 1852 146
rect 2218 143 2252 146
rect 2394 143 2428 146
rect 2570 143 2588 146
rect 2850 143 2868 146
rect 268 133 293 136
rect 290 106 293 133
rect 394 133 404 136
rect 394 116 397 133
rect 418 127 421 135
rect 444 133 493 136
rect 412 124 421 127
rect 498 126 501 135
rect 524 133 549 136
rect 698 133 732 136
rect 770 133 812 136
rect 858 133 868 136
rect 1154 133 1196 136
rect 1338 133 1372 136
rect 1514 133 1540 136
rect 1674 133 1700 136
rect 1842 133 1860 136
rect 1986 133 2028 136
rect 2076 133 2117 136
rect 2260 133 2293 136
rect 2436 133 2469 136
rect 2596 133 2613 136
rect 2740 133 2749 136
rect 2876 133 2901 136
rect 490 123 501 126
rect 564 123 573 126
rect 612 123 645 126
rect 762 123 804 126
rect 842 123 876 126
rect 1092 123 1109 126
rect 1204 123 1221 126
rect 1276 123 1301 126
rect 1452 123 1477 126
rect 1612 123 1637 126
rect 1708 123 1733 126
rect 1772 123 1797 126
rect 1868 123 1877 126
rect 1924 123 1949 126
rect 2084 123 2101 126
rect 2212 123 2221 126
rect 2268 123 2277 126
rect 490 116 493 123
rect 348 113 397 116
rect 444 113 493 116
rect 642 116 645 123
rect 642 113 668 116
rect 692 113 725 116
rect 290 103 340 106
rect 626 103 684 106
rect 14 67 3066 73
rect 38 37 3042 57
rect 14 13 3066 33
<< metal2 >>
rect 2 3033 45 3036
rect 2 6 5 3033
rect 14 13 34 3027
rect 42 3013 45 3033
rect 38 37 58 3003
rect 114 2956 117 3026
rect 106 2953 117 2956
rect 106 2906 109 2953
rect 354 2946 357 2996
rect 130 2923 133 2936
rect 178 2923 181 2946
rect 106 2903 133 2906
rect 130 2646 133 2903
rect 194 2706 197 2926
rect 258 2856 261 2936
rect 290 2933 293 2946
rect 354 2943 365 2946
rect 274 2923 293 2926
rect 330 2923 333 2936
rect 258 2853 269 2856
rect 186 2703 197 2706
rect 130 2643 141 2646
rect 106 2553 109 2606
rect 138 2596 141 2643
rect 130 2593 141 2596
rect 154 2593 157 2616
rect 186 2596 189 2703
rect 202 2696 205 2746
rect 210 2723 213 2766
rect 218 2733 221 2816
rect 266 2776 269 2853
rect 258 2773 269 2776
rect 258 2743 261 2773
rect 202 2693 213 2696
rect 210 2603 213 2693
rect 186 2593 197 2596
rect 66 2236 69 2256
rect 66 2233 77 2236
rect 74 1856 77 2233
rect 66 1853 77 1856
rect 66 1746 69 1853
rect 98 1836 101 2396
rect 130 1843 133 2593
rect 162 2533 165 2556
rect 194 2406 197 2593
rect 226 2566 229 2726
rect 242 2683 245 2736
rect 258 2723 261 2736
rect 282 2713 285 2726
rect 290 2616 293 2923
rect 314 2873 317 2916
rect 362 2896 365 2943
rect 378 2923 381 2946
rect 354 2893 365 2896
rect 306 2763 309 2816
rect 274 2613 297 2616
rect 266 2593 269 2606
rect 226 2563 237 2566
rect 210 2523 213 2536
rect 234 2486 237 2563
rect 226 2483 237 2486
rect 226 2426 229 2483
rect 226 2423 237 2426
rect 186 2403 197 2406
rect 258 2403 261 2566
rect 294 2556 297 2613
rect 294 2553 301 2556
rect 274 2543 285 2546
rect 274 2523 277 2543
rect 282 2533 293 2536
rect 282 2516 285 2526
rect 298 2523 301 2553
rect 306 2533 309 2686
rect 354 2646 357 2893
rect 410 2816 413 2926
rect 410 2813 429 2816
rect 434 2813 437 2876
rect 426 2806 429 2813
rect 410 2793 413 2806
rect 426 2803 437 2806
rect 370 2733 373 2746
rect 378 2683 381 2726
rect 386 2713 389 2736
rect 394 2723 397 2766
rect 434 2753 437 2796
rect 354 2643 365 2646
rect 314 2593 317 2606
rect 330 2553 333 2606
rect 330 2536 333 2546
rect 314 2533 333 2536
rect 346 2526 349 2596
rect 362 2576 365 2643
rect 378 2613 381 2626
rect 402 2603 405 2736
rect 410 2613 413 2636
rect 314 2516 317 2526
rect 282 2513 317 2516
rect 338 2523 349 2526
rect 354 2573 365 2576
rect 266 2443 293 2446
rect 266 2413 269 2443
rect 282 2413 285 2426
rect 290 2416 293 2443
rect 290 2413 301 2416
rect 338 2413 341 2523
rect 266 2403 277 2406
rect 186 2333 189 2403
rect 266 2396 269 2403
rect 234 2393 269 2396
rect 234 2323 237 2393
rect 250 2366 253 2386
rect 250 2363 261 2366
rect 258 2286 261 2363
rect 298 2323 301 2413
rect 354 2406 357 2573
rect 410 2556 413 2576
rect 370 2533 373 2556
rect 406 2553 413 2556
rect 370 2413 373 2516
rect 394 2513 397 2526
rect 406 2496 409 2553
rect 402 2493 409 2496
rect 402 2426 405 2493
rect 402 2423 409 2426
rect 330 2403 357 2406
rect 330 2326 333 2403
rect 354 2346 357 2396
rect 354 2343 373 2346
rect 306 2323 333 2326
rect 354 2323 373 2326
rect 250 2283 261 2286
rect 250 2236 253 2283
rect 242 2233 253 2236
rect 202 2156 205 2176
rect 242 2156 245 2233
rect 274 2186 277 2206
rect 266 2183 277 2186
rect 266 2173 269 2183
rect 162 2153 213 2156
rect 242 2153 253 2156
rect 162 1876 165 2153
rect 210 2133 213 2153
rect 250 2136 253 2153
rect 234 2133 253 2136
rect 234 2086 237 2133
rect 202 2083 237 2086
rect 186 1933 189 2016
rect 202 1976 205 2083
rect 250 2023 253 2126
rect 290 2123 293 2146
rect 306 2126 309 2323
rect 378 2283 381 2336
rect 394 2323 397 2406
rect 406 2306 409 2423
rect 418 2413 421 2746
rect 442 2743 445 2936
rect 466 2933 469 2946
rect 450 2906 453 2926
rect 450 2903 457 2906
rect 454 2836 457 2903
rect 474 2846 477 2936
rect 498 2923 509 2926
rect 522 2916 525 2926
rect 490 2913 525 2916
rect 466 2843 477 2846
rect 454 2833 461 2836
rect 458 2776 461 2833
rect 466 2793 469 2843
rect 458 2773 469 2776
rect 442 2723 445 2736
rect 466 2686 469 2773
rect 506 2756 509 2816
rect 514 2773 525 2776
rect 450 2683 469 2686
rect 426 2563 429 2606
rect 434 2596 437 2616
rect 442 2603 445 2626
rect 450 2613 453 2683
rect 450 2603 461 2606
rect 466 2603 469 2636
rect 474 2596 477 2616
rect 434 2593 477 2596
rect 482 2536 485 2756
rect 506 2753 513 2756
rect 490 2713 493 2726
rect 510 2686 513 2753
rect 522 2696 525 2773
rect 538 2753 541 3016
rect 802 2986 805 3040
rect 782 2983 805 2986
rect 554 2913 557 2936
rect 602 2923 605 2946
rect 626 2923 637 2926
rect 626 2906 629 2923
rect 562 2806 565 2816
rect 546 2803 565 2806
rect 530 2733 533 2746
rect 530 2703 533 2726
rect 538 2723 541 2736
rect 546 2713 549 2736
rect 522 2693 529 2696
rect 506 2683 513 2686
rect 466 2533 485 2536
rect 490 2533 493 2606
rect 506 2603 509 2683
rect 442 2423 445 2436
rect 466 2416 469 2533
rect 482 2506 485 2526
rect 482 2503 493 2506
rect 466 2413 473 2416
rect 418 2316 421 2406
rect 458 2343 461 2396
rect 470 2326 473 2413
rect 490 2376 493 2503
rect 514 2413 517 2616
rect 526 2556 529 2693
rect 554 2666 557 2726
rect 554 2663 565 2666
rect 526 2553 533 2556
rect 522 2513 525 2536
rect 530 2523 533 2553
rect 538 2533 541 2656
rect 546 2593 549 2616
rect 554 2603 557 2636
rect 562 2613 565 2663
rect 570 2616 573 2736
rect 578 2653 581 2806
rect 586 2733 605 2736
rect 618 2733 621 2906
rect 626 2903 633 2906
rect 630 2826 633 2903
rect 626 2823 633 2826
rect 626 2803 629 2823
rect 634 2743 637 2766
rect 602 2703 605 2733
rect 642 2713 645 2936
rect 674 2933 677 2946
rect 658 2776 661 2926
rect 682 2903 685 2936
rect 714 2933 733 2936
rect 714 2926 717 2933
rect 698 2923 717 2926
rect 722 2916 725 2926
rect 690 2913 725 2916
rect 674 2783 677 2806
rect 730 2803 733 2933
rect 738 2896 741 2956
rect 754 2923 757 2936
rect 782 2896 785 2983
rect 826 2966 829 3040
rect 738 2893 749 2896
rect 746 2796 749 2893
rect 778 2893 785 2896
rect 794 2963 829 2966
rect 762 2813 765 2826
rect 778 2796 781 2893
rect 738 2793 749 2796
rect 770 2793 781 2796
rect 650 2773 661 2776
rect 650 2733 653 2773
rect 674 2763 717 2766
rect 738 2763 741 2793
rect 674 2733 677 2763
rect 650 2716 653 2726
rect 658 2723 669 2726
rect 650 2713 677 2716
rect 570 2613 589 2616
rect 626 2613 629 2636
rect 690 2626 693 2736
rect 714 2723 717 2763
rect 770 2736 773 2793
rect 762 2733 773 2736
rect 786 2733 789 2746
rect 682 2623 693 2626
rect 562 2603 573 2606
rect 546 2533 549 2566
rect 466 2323 473 2326
rect 482 2373 493 2376
rect 482 2323 485 2373
rect 490 2353 517 2356
rect 418 2313 429 2316
rect 402 2303 409 2306
rect 322 2253 365 2256
rect 322 2213 325 2253
rect 346 2213 357 2216
rect 362 2213 365 2253
rect 402 2226 405 2303
rect 426 2236 429 2313
rect 418 2233 429 2236
rect 466 2236 469 2323
rect 466 2233 477 2236
rect 402 2223 409 2226
rect 394 2163 397 2206
rect 406 2166 409 2223
rect 418 2213 421 2233
rect 474 2213 477 2233
rect 418 2193 421 2206
rect 434 2203 461 2206
rect 490 2203 493 2353
rect 498 2333 501 2346
rect 514 2333 517 2353
rect 514 2213 517 2326
rect 546 2323 549 2406
rect 562 2403 565 2556
rect 586 2546 589 2613
rect 602 2553 605 2606
rect 682 2576 685 2623
rect 722 2616 725 2726
rect 586 2543 621 2546
rect 594 2423 597 2526
rect 610 2413 613 2536
rect 618 2523 621 2543
rect 626 2533 629 2576
rect 682 2573 693 2576
rect 690 2556 693 2573
rect 698 2563 701 2616
rect 722 2613 733 2616
rect 738 2603 741 2696
rect 762 2626 765 2733
rect 778 2693 781 2726
rect 794 2646 797 2963
rect 906 2956 909 3040
rect 1018 2966 1021 3040
rect 1114 3026 1117 3040
rect 882 2943 885 2956
rect 890 2953 909 2956
rect 1010 2963 1021 2966
rect 1106 3023 1117 3026
rect 802 2886 805 2926
rect 834 2913 837 2926
rect 842 2903 845 2936
rect 858 2913 861 2926
rect 882 2906 885 2926
rect 858 2903 885 2906
rect 802 2883 837 2886
rect 802 2696 805 2766
rect 810 2733 813 2806
rect 818 2783 821 2816
rect 834 2803 837 2883
rect 858 2823 861 2903
rect 866 2803 869 2856
rect 890 2836 893 2953
rect 898 2873 901 2936
rect 930 2853 933 2926
rect 946 2913 949 2936
rect 970 2933 973 2946
rect 890 2833 925 2836
rect 914 2803 917 2826
rect 922 2796 925 2833
rect 946 2823 981 2826
rect 946 2813 949 2823
rect 918 2793 925 2796
rect 834 2763 877 2766
rect 834 2733 837 2763
rect 810 2716 813 2726
rect 818 2723 829 2726
rect 810 2713 837 2716
rect 802 2693 829 2696
rect 794 2643 813 2646
rect 762 2623 805 2626
rect 690 2553 701 2556
rect 698 2533 701 2553
rect 594 2296 597 2326
rect 586 2293 597 2296
rect 406 2163 413 2166
rect 410 2146 413 2163
rect 298 2123 309 2126
rect 234 2013 245 2016
rect 202 1973 213 1976
rect 202 1933 205 1946
rect 138 1873 165 1876
rect 138 1836 141 1873
rect 82 1833 101 1836
rect 130 1833 141 1836
rect 146 1853 189 1856
rect 82 1766 85 1833
rect 98 1793 101 1806
rect 82 1763 93 1766
rect 66 1743 77 1746
rect 74 1496 77 1743
rect 66 1493 77 1496
rect 66 1436 69 1493
rect 90 1476 93 1763
rect 82 1473 93 1476
rect 82 1453 85 1473
rect 66 1433 85 1436
rect 130 1433 133 1833
rect 146 1813 149 1853
rect 170 1813 181 1816
rect 186 1813 189 1853
rect 194 1803 205 1806
rect 154 1523 157 1606
rect 194 1603 197 1626
rect 82 1246 85 1433
rect 138 1366 141 1406
rect 74 1243 85 1246
rect 106 1363 141 1366
rect 74 1176 77 1243
rect 106 1183 109 1363
rect 74 1173 85 1176
rect 82 536 85 1173
rect 138 1166 141 1356
rect 154 1213 157 1226
rect 170 1176 173 1456
rect 186 1393 189 1416
rect 210 1356 213 1973
rect 226 1923 229 1946
rect 250 1873 253 1936
rect 250 1813 253 1866
rect 242 1786 245 1806
rect 234 1783 245 1786
rect 234 1696 237 1783
rect 258 1706 261 2046
rect 298 2026 301 2123
rect 290 2023 301 2026
rect 322 2026 325 2136
rect 370 2123 373 2146
rect 410 2143 421 2146
rect 394 2133 413 2136
rect 322 2023 333 2026
rect 290 1926 293 2023
rect 314 2006 317 2016
rect 306 2003 317 2006
rect 266 1906 269 1926
rect 290 1923 301 1926
rect 314 1923 317 2003
rect 330 1966 333 2023
rect 394 2013 397 2133
rect 418 2126 421 2143
rect 410 2123 421 2126
rect 402 2013 405 2036
rect 322 1963 333 1966
rect 266 1903 277 1906
rect 274 1846 277 1903
rect 298 1893 301 1923
rect 322 1856 325 1963
rect 370 1956 373 2006
rect 362 1953 373 1956
rect 330 1933 333 1946
rect 330 1913 349 1916
rect 346 1856 349 1913
rect 362 1866 365 1953
rect 386 1923 389 1936
rect 362 1863 369 1866
rect 266 1843 277 1846
rect 298 1853 325 1856
rect 338 1853 349 1856
rect 266 1823 269 1843
rect 282 1803 285 1826
rect 298 1766 301 1853
rect 322 1813 325 1826
rect 338 1776 341 1853
rect 366 1806 369 1863
rect 378 1813 381 1876
rect 410 1826 413 2123
rect 418 2013 421 2026
rect 426 2023 429 2126
rect 418 1923 421 2006
rect 434 1913 437 2126
rect 442 2116 445 2126
rect 442 2113 453 2116
rect 442 2033 445 2106
rect 450 2083 453 2113
rect 458 1836 461 2203
rect 466 2133 469 2146
rect 474 2113 477 2166
rect 570 2136 573 2216
rect 586 2206 589 2293
rect 618 2286 621 2356
rect 642 2323 645 2336
rect 482 2093 485 2136
rect 522 2106 525 2136
rect 562 2133 573 2136
rect 578 2203 589 2206
rect 602 2283 621 2286
rect 602 2203 605 2283
rect 626 2213 629 2286
rect 650 2256 653 2436
rect 674 2413 677 2426
rect 682 2393 685 2446
rect 730 2413 733 2576
rect 754 2573 757 2606
rect 770 2583 773 2616
rect 778 2613 789 2616
rect 778 2566 781 2606
rect 786 2603 797 2606
rect 746 2563 781 2566
rect 746 2523 749 2563
rect 794 2513 797 2586
rect 794 2413 797 2426
rect 714 2393 717 2406
rect 738 2373 741 2396
rect 778 2393 797 2396
rect 642 2253 653 2256
rect 514 2103 525 2106
rect 514 2036 517 2103
rect 498 2033 517 2036
rect 482 2023 509 2026
rect 466 1926 469 1946
rect 482 1936 485 2023
rect 514 2016 517 2026
rect 490 2013 517 2016
rect 482 1933 489 1936
rect 466 1923 477 1926
rect 458 1833 465 1836
rect 402 1823 413 1826
rect 366 1803 373 1806
rect 338 1773 349 1776
rect 274 1763 301 1766
rect 274 1733 277 1763
rect 322 1723 325 1746
rect 346 1736 349 1773
rect 342 1733 349 1736
rect 258 1703 269 1706
rect 234 1693 245 1696
rect 218 1613 221 1626
rect 218 1513 221 1526
rect 242 1523 245 1693
rect 258 1603 261 1616
rect 258 1533 261 1546
rect 130 1163 141 1166
rect 154 1173 173 1176
rect 194 1353 213 1356
rect 130 716 133 1163
rect 154 723 157 1173
rect 194 1026 197 1353
rect 226 1296 229 1436
rect 234 1413 237 1506
rect 250 1456 253 1526
rect 266 1516 269 1703
rect 342 1686 345 1733
rect 338 1683 345 1686
rect 338 1626 341 1683
rect 306 1623 341 1626
rect 282 1603 285 1616
rect 306 1556 309 1623
rect 346 1613 349 1626
rect 354 1606 357 1726
rect 370 1723 373 1803
rect 402 1766 405 1823
rect 450 1816 453 1826
rect 418 1793 421 1816
rect 434 1813 453 1816
rect 402 1763 413 1766
rect 394 1733 397 1746
rect 402 1676 405 1696
rect 386 1673 405 1676
rect 338 1603 357 1606
rect 362 1566 365 1626
rect 354 1563 365 1566
rect 306 1553 325 1556
rect 282 1543 301 1546
rect 282 1536 285 1543
rect 274 1533 285 1536
rect 266 1513 277 1516
rect 246 1453 253 1456
rect 246 1356 249 1453
rect 246 1353 253 1356
rect 210 1293 229 1296
rect 210 1206 213 1293
rect 250 1286 253 1353
rect 226 1283 253 1286
rect 226 1213 229 1283
rect 250 1223 253 1246
rect 234 1213 245 1216
rect 258 1213 261 1446
rect 266 1313 269 1326
rect 210 1203 221 1206
rect 218 1036 221 1203
rect 234 1133 237 1213
rect 266 1186 269 1296
rect 274 1276 277 1513
rect 282 1503 285 1526
rect 290 1473 293 1536
rect 298 1533 301 1543
rect 298 1336 301 1526
rect 322 1446 325 1553
rect 354 1523 357 1563
rect 386 1556 389 1673
rect 410 1656 413 1763
rect 426 1756 429 1806
rect 418 1733 421 1756
rect 426 1753 441 1756
rect 426 1723 429 1746
rect 402 1653 413 1656
rect 402 1576 405 1653
rect 418 1633 421 1716
rect 402 1573 413 1576
rect 386 1553 405 1556
rect 386 1516 389 1536
rect 402 1523 405 1553
rect 290 1333 301 1336
rect 306 1443 325 1446
rect 378 1513 389 1516
rect 306 1336 309 1443
rect 378 1426 381 1513
rect 410 1506 413 1573
rect 418 1523 421 1626
rect 426 1613 429 1676
rect 438 1636 441 1753
rect 438 1633 445 1636
rect 442 1613 445 1633
rect 450 1623 453 1813
rect 462 1616 465 1833
rect 474 1803 477 1923
rect 486 1886 489 1933
rect 506 1923 509 1996
rect 482 1883 489 1886
rect 482 1863 485 1883
rect 506 1876 509 1916
rect 490 1803 493 1816
rect 482 1793 493 1796
rect 474 1643 477 1736
rect 490 1693 493 1793
rect 498 1733 501 1876
rect 506 1873 517 1876
rect 514 1686 517 1873
rect 538 1823 541 2116
rect 562 2023 565 2036
rect 546 2013 573 2016
rect 578 2003 581 2203
rect 642 2176 645 2253
rect 698 2226 701 2326
rect 722 2296 725 2336
rect 674 2223 701 2226
rect 714 2293 725 2296
rect 714 2226 717 2293
rect 746 2266 749 2326
rect 802 2323 805 2623
rect 810 2506 813 2643
rect 826 2626 829 2693
rect 818 2623 829 2626
rect 818 2583 821 2623
rect 826 2573 829 2606
rect 850 2576 853 2736
rect 874 2723 877 2763
rect 834 2573 853 2576
rect 834 2566 837 2573
rect 826 2563 837 2566
rect 826 2533 829 2563
rect 850 2516 853 2566
rect 858 2553 861 2616
rect 874 2613 877 2716
rect 882 2606 885 2776
rect 890 2613 893 2726
rect 918 2686 921 2793
rect 930 2763 933 2806
rect 946 2773 949 2806
rect 954 2793 957 2816
rect 962 2796 965 2806
rect 970 2803 973 2816
rect 978 2803 981 2823
rect 994 2796 997 2926
rect 1010 2896 1013 2963
rect 1066 2933 1069 2946
rect 1042 2923 1053 2926
rect 1010 2893 1021 2896
rect 1010 2803 1013 2876
rect 1018 2866 1021 2893
rect 1042 2873 1045 2923
rect 1018 2863 1053 2866
rect 962 2793 997 2796
rect 1018 2793 1021 2816
rect 946 2733 949 2756
rect 914 2683 921 2686
rect 898 2606 901 2636
rect 914 2606 917 2683
rect 930 2633 933 2726
rect 954 2706 957 2726
rect 962 2713 965 2736
rect 970 2723 973 2786
rect 978 2733 981 2776
rect 1034 2763 1037 2806
rect 978 2723 989 2726
rect 978 2706 981 2723
rect 954 2703 981 2706
rect 986 2656 989 2723
rect 994 2693 997 2736
rect 1018 2666 1021 2736
rect 1042 2713 1045 2726
rect 1018 2663 1037 2666
rect 986 2653 1017 2656
rect 994 2613 997 2636
rect 866 2523 869 2606
rect 874 2603 885 2606
rect 890 2603 901 2606
rect 906 2603 917 2606
rect 850 2513 869 2516
rect 810 2503 821 2506
rect 818 2476 821 2503
rect 818 2473 829 2476
rect 826 2376 829 2473
rect 866 2413 869 2513
rect 906 2436 909 2603
rect 922 2523 925 2556
rect 938 2516 941 2546
rect 946 2533 949 2606
rect 1014 2556 1017 2653
rect 1034 2606 1037 2663
rect 1026 2603 1037 2606
rect 970 2523 973 2556
rect 1014 2553 1021 2556
rect 978 2516 981 2546
rect 898 2433 909 2436
rect 850 2403 861 2406
rect 818 2373 829 2376
rect 818 2356 821 2373
rect 814 2353 821 2356
rect 814 2306 817 2353
rect 834 2333 837 2356
rect 858 2323 861 2403
rect 874 2373 877 2396
rect 898 2386 901 2433
rect 914 2403 917 2426
rect 930 2413 933 2516
rect 938 2513 981 2516
rect 938 2496 941 2513
rect 938 2493 949 2496
rect 946 2436 949 2493
rect 1010 2473 1013 2536
rect 1018 2526 1021 2553
rect 1026 2533 1029 2603
rect 1034 2543 1037 2586
rect 1050 2546 1053 2863
rect 1074 2766 1077 2886
rect 1090 2836 1093 2926
rect 1106 2886 1109 3023
rect 1130 2966 1133 3040
rect 1450 2993 1453 3040
rect 1130 2963 1137 2966
rect 1134 2886 1137 2963
rect 1146 2913 1149 2926
rect 1106 2883 1117 2886
rect 1082 2833 1093 2836
rect 1082 2803 1085 2833
rect 1114 2816 1117 2883
rect 1130 2883 1137 2886
rect 1162 2883 1165 2926
rect 1090 2793 1093 2816
rect 1114 2813 1121 2816
rect 1074 2763 1085 2766
rect 1066 2736 1069 2756
rect 1062 2733 1069 2736
rect 1062 2686 1065 2733
rect 1082 2723 1085 2763
rect 1098 2736 1101 2806
rect 1090 2733 1101 2736
rect 1106 2733 1109 2806
rect 1118 2756 1121 2813
rect 1114 2753 1121 2756
rect 1130 2756 1133 2883
rect 1282 2856 1285 2946
rect 1266 2853 1285 2856
rect 1298 2873 1309 2876
rect 1154 2833 1189 2836
rect 1154 2813 1157 2833
rect 1162 2803 1165 2826
rect 1170 2793 1173 2816
rect 1130 2753 1157 2756
rect 1114 2733 1117 2753
rect 1130 2743 1141 2746
rect 1122 2733 1133 2736
rect 1138 2733 1141 2743
rect 1146 2733 1149 2746
rect 1062 2683 1069 2686
rect 1066 2606 1069 2683
rect 1090 2666 1093 2733
rect 1098 2693 1101 2726
rect 1114 2713 1117 2726
rect 1122 2723 1133 2726
rect 1146 2713 1149 2726
rect 1154 2706 1157 2753
rect 1170 2733 1173 2786
rect 1178 2773 1181 2806
rect 1186 2776 1189 2833
rect 1250 2813 1253 2826
rect 1202 2803 1213 2806
rect 1226 2783 1229 2806
rect 1186 2773 1241 2776
rect 1194 2723 1197 2736
rect 1238 2716 1241 2773
rect 1250 2723 1253 2746
rect 1266 2733 1269 2853
rect 1298 2826 1301 2873
rect 1294 2823 1301 2826
rect 1138 2703 1157 2706
rect 1090 2663 1109 2666
rect 1066 2603 1077 2606
rect 1074 2573 1077 2603
rect 1046 2543 1053 2546
rect 1018 2523 1029 2526
rect 1034 2513 1037 2536
rect 1046 2496 1049 2543
rect 1042 2493 1049 2496
rect 938 2433 949 2436
rect 1042 2436 1045 2493
rect 1042 2433 1053 2436
rect 914 2386 917 2396
rect 938 2386 941 2433
rect 954 2403 957 2416
rect 994 2413 997 2426
rect 898 2383 909 2386
rect 914 2383 941 2386
rect 882 2306 885 2366
rect 906 2326 909 2383
rect 922 2333 925 2383
rect 946 2343 949 2396
rect 970 2363 973 2406
rect 1050 2396 1053 2433
rect 1042 2393 1053 2396
rect 814 2303 821 2306
rect 730 2263 749 2266
rect 714 2223 725 2226
rect 642 2173 653 2176
rect 602 2123 637 2126
rect 594 1933 597 2066
rect 602 2036 605 2116
rect 618 2083 621 2116
rect 602 2033 621 2036
rect 602 2013 605 2033
rect 554 1846 557 1926
rect 586 1873 589 1926
rect 618 1923 621 2033
rect 634 2013 637 2123
rect 650 2043 653 2173
rect 674 2146 677 2223
rect 674 2143 681 2146
rect 666 2076 669 2136
rect 678 2086 681 2143
rect 658 2073 669 2076
rect 674 2083 681 2086
rect 650 1996 653 2026
rect 642 1993 653 1996
rect 642 1936 645 1993
rect 658 1963 661 2073
rect 674 2066 677 2083
rect 666 2063 677 2066
rect 666 2046 669 2063
rect 666 2043 673 2046
rect 670 1946 673 2043
rect 690 2036 693 2216
rect 706 2126 709 2206
rect 722 2186 725 2223
rect 730 2213 733 2263
rect 794 2213 797 2226
rect 818 2216 821 2303
rect 874 2303 885 2306
rect 898 2323 917 2326
rect 874 2226 877 2303
rect 818 2213 829 2216
rect 834 2213 837 2226
rect 874 2223 885 2226
rect 746 2186 749 2206
rect 722 2183 749 2186
rect 746 2176 749 2183
rect 770 2176 773 2186
rect 746 2173 773 2176
rect 722 2133 741 2136
rect 738 2126 741 2133
rect 706 2123 717 2126
rect 698 2093 701 2116
rect 714 2113 717 2123
rect 730 2073 733 2126
rect 738 2123 749 2126
rect 738 2113 749 2116
rect 754 2096 757 2136
rect 746 2093 757 2096
rect 626 1933 645 1936
rect 666 1943 673 1946
rect 682 2033 693 2036
rect 626 1906 629 1933
rect 666 1926 669 1943
rect 618 1903 629 1906
rect 554 1843 581 1846
rect 546 1823 573 1826
rect 538 1803 541 1816
rect 546 1813 549 1823
rect 554 1766 557 1816
rect 562 1813 573 1816
rect 578 1803 581 1843
rect 618 1826 621 1903
rect 618 1823 629 1826
rect 618 1783 621 1806
rect 506 1683 517 1686
rect 546 1763 557 1766
rect 458 1613 465 1616
rect 410 1503 421 1506
rect 314 1423 341 1426
rect 378 1423 389 1426
rect 314 1413 317 1423
rect 322 1403 325 1416
rect 306 1333 317 1336
rect 330 1333 333 1423
rect 338 1393 341 1406
rect 290 1293 293 1333
rect 298 1323 309 1326
rect 274 1273 281 1276
rect 258 1183 269 1186
rect 258 1126 261 1183
rect 278 1176 281 1273
rect 314 1243 317 1333
rect 346 1313 349 1326
rect 290 1213 293 1226
rect 298 1203 301 1226
rect 370 1213 373 1226
rect 386 1216 389 1423
rect 402 1413 405 1476
rect 418 1406 421 1503
rect 410 1403 421 1406
rect 434 1403 437 1606
rect 450 1516 453 1536
rect 446 1513 453 1516
rect 446 1426 449 1513
rect 446 1423 453 1426
rect 410 1346 413 1403
rect 450 1373 453 1423
rect 402 1343 413 1346
rect 402 1236 405 1343
rect 402 1233 413 1236
rect 386 1213 405 1216
rect 322 1183 325 1206
rect 274 1173 281 1176
rect 258 1123 269 1126
rect 266 1103 269 1123
rect 218 1033 253 1036
rect 194 1023 213 1026
rect 130 713 141 716
rect 66 533 85 536
rect 66 513 69 533
rect 66 416 69 436
rect 66 413 85 416
rect 82 6 85 413
rect 138 13 141 713
rect 210 623 213 1023
rect 250 856 253 1033
rect 242 853 253 856
rect 242 776 245 853
rect 234 773 245 776
rect 234 716 237 773
rect 274 766 277 1173
rect 282 1013 285 1126
rect 322 1013 333 1016
rect 370 976 373 1186
rect 394 1123 397 1156
rect 394 993 397 1016
rect 354 973 373 976
rect 322 933 325 956
rect 290 813 293 916
rect 354 856 357 973
rect 378 866 381 916
rect 394 903 397 936
rect 410 916 413 1233
rect 418 1203 421 1336
rect 426 1176 429 1306
rect 434 1183 437 1336
rect 458 1303 461 1613
rect 490 1596 493 1626
rect 482 1593 493 1596
rect 498 1596 501 1606
rect 506 1603 509 1683
rect 546 1666 549 1763
rect 562 1673 565 1736
rect 570 1733 573 1776
rect 626 1746 629 1823
rect 642 1813 645 1926
rect 650 1913 653 1926
rect 658 1923 669 1926
rect 674 1916 677 1926
rect 666 1913 677 1916
rect 666 1816 669 1913
rect 658 1813 669 1816
rect 586 1743 629 1746
rect 634 1803 645 1806
rect 546 1663 557 1666
rect 530 1596 533 1606
rect 498 1593 533 1596
rect 482 1536 485 1593
rect 482 1533 493 1536
rect 466 1513 485 1516
rect 466 1496 469 1513
rect 466 1493 473 1496
rect 470 1426 473 1493
rect 490 1473 493 1533
rect 506 1506 509 1546
rect 530 1523 533 1536
rect 538 1523 541 1626
rect 554 1603 557 1663
rect 586 1593 589 1743
rect 610 1706 613 1736
rect 634 1716 637 1803
rect 658 1746 661 1813
rect 674 1756 677 1806
rect 682 1773 685 2033
rect 698 1993 701 2006
rect 722 1933 725 2016
rect 746 2013 749 2093
rect 762 1933 765 2086
rect 698 1906 701 1926
rect 754 1906 757 1926
rect 698 1903 709 1906
rect 706 1826 709 1903
rect 746 1903 757 1906
rect 746 1846 749 1903
rect 746 1843 757 1846
rect 674 1753 681 1756
rect 658 1743 669 1746
rect 650 1716 653 1726
rect 666 1716 669 1743
rect 618 1713 629 1716
rect 610 1703 621 1706
rect 618 1636 621 1703
rect 614 1633 621 1636
rect 602 1546 605 1606
rect 614 1556 617 1633
rect 626 1566 629 1713
rect 634 1713 645 1716
rect 650 1713 669 1716
rect 634 1583 637 1713
rect 626 1563 633 1566
rect 614 1553 621 1556
rect 546 1533 549 1546
rect 594 1543 605 1546
rect 594 1526 597 1543
rect 506 1503 517 1506
rect 514 1436 517 1503
rect 578 1473 581 1526
rect 590 1523 597 1526
rect 602 1523 605 1536
rect 618 1533 621 1553
rect 506 1433 517 1436
rect 590 1436 593 1523
rect 590 1433 597 1436
rect 466 1423 473 1426
rect 466 1333 469 1423
rect 498 1416 501 1426
rect 482 1413 501 1416
rect 506 1413 509 1433
rect 594 1413 597 1433
rect 482 1336 485 1413
rect 602 1406 605 1516
rect 554 1386 557 1406
rect 546 1383 557 1386
rect 586 1403 605 1406
rect 474 1333 485 1336
rect 474 1316 477 1333
rect 470 1313 477 1316
rect 470 1246 473 1313
rect 482 1266 485 1326
rect 514 1323 517 1376
rect 546 1323 549 1383
rect 586 1336 589 1403
rect 618 1383 621 1526
rect 630 1496 633 1563
rect 626 1493 633 1496
rect 578 1333 589 1336
rect 578 1276 581 1333
rect 594 1286 597 1326
rect 626 1323 629 1493
rect 642 1486 645 1636
rect 650 1626 653 1706
rect 658 1633 661 1656
rect 650 1623 661 1626
rect 650 1603 653 1616
rect 658 1586 661 1623
rect 666 1606 669 1713
rect 678 1696 681 1753
rect 690 1713 693 1826
rect 698 1823 709 1826
rect 698 1803 701 1823
rect 714 1733 717 1766
rect 678 1693 685 1696
rect 682 1616 685 1693
rect 738 1686 741 1816
rect 746 1803 749 1826
rect 754 1743 757 1843
rect 762 1803 765 1866
rect 770 1763 773 2173
rect 794 2133 797 2146
rect 826 2133 829 2166
rect 778 2106 781 2126
rect 802 2123 813 2126
rect 778 2103 789 2106
rect 802 2103 805 2123
rect 842 2116 845 2206
rect 874 2186 877 2206
rect 870 2183 877 2186
rect 810 2113 853 2116
rect 786 2036 789 2103
rect 778 2033 789 2036
rect 778 2013 781 2033
rect 810 2013 813 2113
rect 802 2003 813 2006
rect 778 1976 781 1996
rect 778 1973 785 1976
rect 782 1836 785 1973
rect 802 1956 805 2003
rect 802 1953 809 1956
rect 794 1873 797 1926
rect 806 1886 809 1953
rect 818 1896 821 2096
rect 858 2013 861 2136
rect 870 2016 873 2183
rect 870 2013 877 2016
rect 834 1993 837 2006
rect 826 1933 829 1946
rect 874 1933 877 2013
rect 882 1976 885 2223
rect 898 2203 901 2323
rect 1034 2306 1037 2326
rect 1026 2303 1037 2306
rect 906 2196 909 2216
rect 922 2206 925 2216
rect 914 2203 925 2206
rect 898 2193 909 2196
rect 898 2133 901 2193
rect 930 2163 933 2216
rect 938 2193 941 2206
rect 922 2133 925 2146
rect 898 2106 901 2126
rect 946 2116 949 2276
rect 1026 2246 1029 2303
rect 1026 2243 1037 2246
rect 994 2213 1013 2216
rect 962 2126 965 2206
rect 1010 2193 1013 2206
rect 962 2123 1013 2126
rect 938 2113 949 2116
rect 898 2103 909 2106
rect 906 2046 909 2103
rect 898 2043 909 2046
rect 938 2046 941 2113
rect 938 2043 949 2046
rect 898 2026 901 2043
rect 898 2023 925 2026
rect 914 2003 917 2016
rect 946 2006 949 2043
rect 954 2036 957 2116
rect 962 2113 981 2116
rect 962 2103 965 2113
rect 970 2046 973 2106
rect 986 2093 989 2106
rect 970 2043 981 2046
rect 954 2033 965 2036
rect 954 2013 957 2026
rect 962 2013 965 2033
rect 930 2003 949 2006
rect 882 1973 909 1976
rect 834 1913 837 1926
rect 818 1893 829 1896
rect 806 1883 813 1886
rect 778 1833 785 1836
rect 762 1713 765 1726
rect 722 1683 741 1686
rect 682 1613 693 1616
rect 666 1603 677 1606
rect 658 1583 669 1586
rect 642 1483 649 1486
rect 634 1333 637 1476
rect 646 1396 649 1483
rect 666 1456 669 1583
rect 690 1523 693 1613
rect 706 1596 709 1626
rect 722 1613 725 1683
rect 738 1616 741 1626
rect 730 1613 741 1616
rect 746 1616 749 1646
rect 746 1613 757 1616
rect 730 1596 733 1613
rect 706 1593 733 1596
rect 746 1593 749 1606
rect 658 1453 669 1456
rect 658 1413 661 1453
rect 690 1413 693 1516
rect 706 1443 709 1526
rect 738 1513 741 1586
rect 754 1573 757 1613
rect 778 1606 781 1833
rect 786 1723 789 1816
rect 802 1793 805 1816
rect 810 1803 813 1883
rect 826 1796 829 1893
rect 818 1793 829 1796
rect 818 1736 821 1793
rect 794 1723 797 1736
rect 802 1733 813 1736
rect 818 1733 829 1736
rect 802 1713 805 1726
rect 794 1613 797 1676
rect 810 1613 813 1733
rect 826 1606 829 1733
rect 770 1556 773 1606
rect 778 1603 797 1606
rect 762 1553 773 1556
rect 762 1506 765 1553
rect 762 1503 773 1506
rect 738 1413 741 1426
rect 754 1413 757 1426
rect 770 1423 773 1503
rect 794 1446 797 1603
rect 810 1583 813 1606
rect 826 1603 837 1606
rect 826 1523 829 1596
rect 786 1443 797 1446
rect 834 1443 837 1603
rect 666 1403 685 1406
rect 646 1393 653 1396
rect 650 1346 653 1393
rect 642 1343 653 1346
rect 642 1323 645 1343
rect 682 1326 685 1403
rect 722 1333 733 1336
rect 666 1306 669 1326
rect 682 1323 725 1326
rect 650 1303 669 1306
rect 594 1283 605 1286
rect 578 1273 589 1276
rect 482 1263 525 1266
rect 470 1243 477 1246
rect 442 1203 445 1216
rect 450 1203 453 1226
rect 466 1216 469 1226
rect 458 1213 469 1216
rect 426 1173 453 1176
rect 450 1006 453 1173
rect 466 1013 469 1206
rect 474 1203 477 1243
rect 482 1203 485 1216
rect 522 1203 525 1263
rect 530 1213 533 1226
rect 546 1203 549 1216
rect 450 1003 461 1006
rect 410 913 429 916
rect 378 863 385 866
rect 338 853 357 856
rect 314 813 325 816
rect 338 776 341 853
rect 354 793 357 806
rect 382 796 385 863
rect 418 856 421 906
rect 434 893 437 936
rect 458 933 461 1003
rect 482 923 485 1026
rect 490 996 493 1186
rect 530 1133 533 1176
rect 546 1133 549 1156
rect 562 1133 565 1206
rect 586 1203 589 1273
rect 514 1013 517 1126
rect 530 1013 533 1126
rect 546 1123 557 1126
rect 594 1123 597 1216
rect 602 1203 605 1283
rect 546 1013 549 1123
rect 490 993 501 996
rect 538 993 541 1006
rect 554 1003 557 1016
rect 562 1013 565 1036
rect 498 916 501 993
rect 538 943 557 946
rect 586 943 589 1036
rect 602 1003 605 1156
rect 610 1123 613 1216
rect 618 1116 621 1226
rect 626 1196 629 1216
rect 626 1193 637 1196
rect 634 1146 637 1193
rect 626 1143 637 1146
rect 626 1123 629 1143
rect 650 1136 653 1303
rect 674 1286 677 1316
rect 682 1296 685 1316
rect 682 1293 693 1296
rect 666 1283 677 1286
rect 666 1226 669 1283
rect 690 1246 693 1293
rect 682 1243 693 1246
rect 666 1223 677 1226
rect 674 1203 677 1223
rect 682 1156 685 1243
rect 690 1203 693 1216
rect 698 1173 701 1216
rect 682 1153 693 1156
rect 650 1133 661 1136
rect 618 1113 637 1116
rect 658 1036 661 1133
rect 682 1126 685 1146
rect 674 1123 685 1126
rect 658 1033 669 1036
rect 610 1023 621 1026
rect 538 933 541 943
rect 642 933 645 946
rect 490 913 501 916
rect 418 853 437 856
rect 378 793 385 796
rect 338 773 357 776
rect 274 763 301 766
rect 250 753 269 756
rect 250 733 253 753
rect 266 746 269 753
rect 258 723 261 746
rect 266 743 293 746
rect 234 713 245 716
rect 242 476 245 713
rect 234 473 245 476
rect 234 403 237 473
rect 266 413 269 743
rect 274 733 293 736
rect 274 613 277 733
rect 298 666 301 763
rect 290 663 301 666
rect 290 596 293 663
rect 354 646 357 773
rect 378 676 381 793
rect 394 733 397 816
rect 434 813 437 853
rect 450 793 453 806
rect 402 743 405 756
rect 450 723 453 736
rect 474 733 477 816
rect 490 726 493 913
rect 530 813 533 896
rect 618 893 621 926
rect 546 793 549 806
rect 498 743 509 746
rect 514 743 517 756
rect 578 733 581 816
rect 626 813 629 926
rect 658 923 661 1016
rect 666 953 669 1033
rect 674 1023 677 1123
rect 690 1116 693 1153
rect 706 1146 709 1226
rect 706 1143 717 1146
rect 682 1113 693 1116
rect 682 1033 685 1113
rect 690 1096 693 1106
rect 698 1103 701 1116
rect 690 1093 701 1096
rect 698 1056 701 1093
rect 706 1073 709 1136
rect 714 1106 717 1143
rect 722 1123 725 1323
rect 730 1313 733 1326
rect 738 1323 741 1406
rect 746 1393 749 1406
rect 778 1403 781 1416
rect 746 1203 749 1326
rect 762 1313 765 1336
rect 786 1323 789 1443
rect 794 1393 797 1436
rect 794 1316 797 1326
rect 810 1323 813 1336
rect 826 1333 829 1406
rect 834 1336 837 1426
rect 842 1346 845 1916
rect 874 1813 877 1826
rect 858 1733 861 1786
rect 866 1756 869 1806
rect 882 1803 885 1966
rect 906 1826 909 1973
rect 922 1913 925 1946
rect 930 1923 933 2003
rect 938 1916 941 1996
rect 954 1946 957 2006
rect 930 1913 941 1916
rect 946 1943 957 1946
rect 906 1823 917 1826
rect 914 1806 917 1823
rect 890 1793 893 1806
rect 906 1803 917 1806
rect 906 1756 909 1803
rect 866 1753 885 1756
rect 906 1753 917 1756
rect 866 1723 869 1746
rect 858 1533 861 1616
rect 866 1613 869 1646
rect 850 1393 853 1416
rect 874 1366 877 1736
rect 882 1723 885 1753
rect 898 1663 901 1736
rect 914 1706 917 1753
rect 922 1723 925 1806
rect 930 1733 933 1913
rect 946 1836 949 1943
rect 978 1936 981 2043
rect 1002 2016 1005 2116
rect 1018 2083 1021 2206
rect 1026 2113 1029 2226
rect 1034 2196 1037 2243
rect 1042 2203 1045 2393
rect 1058 2336 1061 2536
rect 1082 2523 1085 2616
rect 1090 2603 1093 2636
rect 1098 2613 1101 2656
rect 1106 2603 1109 2663
rect 1114 2586 1117 2596
rect 1106 2583 1117 2586
rect 1138 2556 1141 2703
rect 1138 2553 1157 2556
rect 1098 2533 1101 2546
rect 1074 2363 1077 2406
rect 1098 2403 1101 2416
rect 1114 2363 1117 2536
rect 1138 2456 1141 2553
rect 1146 2523 1149 2546
rect 1162 2536 1165 2706
rect 1194 2613 1197 2716
rect 1238 2713 1245 2716
rect 1242 2613 1245 2713
rect 1294 2686 1297 2823
rect 1306 2803 1309 2816
rect 1314 2796 1317 2976
rect 1386 2933 1389 2946
rect 1330 2893 1333 2926
rect 1338 2826 1341 2846
rect 1266 2683 1297 2686
rect 1306 2793 1317 2796
rect 1330 2823 1341 2826
rect 1186 2586 1189 2606
rect 1158 2533 1165 2536
rect 1182 2583 1189 2586
rect 1158 2486 1161 2533
rect 1182 2516 1185 2583
rect 1202 2573 1205 2596
rect 1194 2523 1197 2556
rect 1182 2513 1189 2516
rect 1186 2493 1189 2513
rect 1210 2486 1213 2536
rect 1234 2513 1237 2526
rect 1158 2483 1165 2486
rect 1138 2453 1149 2456
rect 1146 2376 1149 2453
rect 1130 2373 1149 2376
rect 1058 2333 1077 2336
rect 1050 2323 1061 2326
rect 1050 2226 1053 2323
rect 1058 2303 1061 2316
rect 1066 2233 1069 2306
rect 1050 2223 1061 2226
rect 1074 2216 1077 2333
rect 1082 2303 1085 2336
rect 1090 2296 1093 2316
rect 1122 2306 1125 2326
rect 1114 2303 1125 2306
rect 1090 2293 1101 2296
rect 1058 2213 1077 2216
rect 1034 2193 1045 2196
rect 1042 2123 1045 2193
rect 1058 2106 1061 2213
rect 1098 2206 1101 2293
rect 1114 2236 1117 2303
rect 1114 2233 1125 2236
rect 1130 2233 1133 2373
rect 1162 2346 1165 2483
rect 1186 2483 1213 2486
rect 1186 2363 1189 2483
rect 1210 2413 1213 2476
rect 1250 2456 1253 2616
rect 1266 2576 1269 2683
rect 1306 2676 1309 2793
rect 1330 2776 1333 2823
rect 1346 2803 1349 2916
rect 1370 2913 1373 2926
rect 1386 2836 1389 2926
rect 1382 2833 1389 2836
rect 1330 2773 1341 2776
rect 1354 2773 1357 2816
rect 1370 2813 1373 2826
rect 1382 2786 1385 2833
rect 1394 2796 1397 2826
rect 1402 2803 1405 2896
rect 1434 2886 1437 2926
rect 1434 2883 1461 2886
rect 1394 2793 1405 2796
rect 1382 2783 1389 2786
rect 1338 2756 1341 2773
rect 1338 2753 1349 2756
rect 1282 2673 1309 2676
rect 1266 2573 1277 2576
rect 1274 2536 1277 2573
rect 1282 2556 1285 2673
rect 1314 2616 1317 2726
rect 1346 2686 1349 2753
rect 1370 2706 1373 2726
rect 1338 2683 1349 2686
rect 1362 2703 1373 2706
rect 1290 2566 1293 2606
rect 1298 2603 1301 2616
rect 1314 2613 1325 2616
rect 1322 2603 1325 2613
rect 1338 2576 1341 2683
rect 1362 2656 1365 2703
rect 1362 2653 1373 2656
rect 1354 2623 1357 2636
rect 1346 2613 1365 2616
rect 1370 2613 1373 2653
rect 1378 2613 1381 2726
rect 1386 2706 1389 2783
rect 1394 2723 1397 2736
rect 1402 2723 1405 2793
rect 1426 2736 1429 2826
rect 1442 2793 1445 2806
rect 1434 2736 1437 2746
rect 1450 2736 1453 2836
rect 1458 2816 1461 2883
rect 1466 2843 1469 3040
rect 1482 2936 1485 3040
rect 1506 2996 1509 3040
rect 1522 3023 1525 3040
rect 1506 2993 1513 2996
rect 1478 2933 1485 2936
rect 1478 2886 1481 2933
rect 1474 2883 1481 2886
rect 1474 2833 1477 2883
rect 1490 2876 1493 2926
rect 1482 2873 1493 2876
rect 1458 2813 1469 2816
rect 1466 2803 1469 2813
rect 1426 2733 1437 2736
rect 1410 2723 1421 2726
rect 1386 2703 1397 2706
rect 1346 2593 1349 2613
rect 1394 2606 1397 2703
rect 1410 2653 1413 2723
rect 1426 2713 1429 2726
rect 1426 2613 1429 2636
rect 1338 2573 1345 2576
rect 1290 2563 1333 2566
rect 1282 2553 1293 2556
rect 1274 2533 1281 2536
rect 1278 2486 1281 2533
rect 1274 2483 1281 2486
rect 1250 2453 1261 2456
rect 1258 2376 1261 2453
rect 1250 2373 1261 2376
rect 1162 2343 1181 2346
rect 1154 2323 1173 2326
rect 1162 2273 1165 2316
rect 1138 2233 1157 2236
rect 1170 2233 1173 2323
rect 1178 2303 1181 2343
rect 1250 2323 1253 2373
rect 1274 2356 1277 2483
rect 1290 2463 1293 2553
rect 1306 2456 1309 2536
rect 1330 2523 1333 2563
rect 1342 2496 1345 2573
rect 1298 2453 1309 2456
rect 1298 2363 1301 2453
rect 1322 2413 1325 2496
rect 1338 2493 1345 2496
rect 1338 2473 1341 2493
rect 1354 2466 1357 2606
rect 1386 2603 1397 2606
rect 1378 2536 1381 2556
rect 1374 2533 1381 2536
rect 1374 2476 1377 2533
rect 1386 2483 1389 2603
rect 1418 2583 1421 2606
rect 1426 2576 1429 2606
rect 1434 2593 1437 2733
rect 1446 2733 1453 2736
rect 1446 2646 1449 2733
rect 1442 2643 1449 2646
rect 1426 2573 1433 2576
rect 1402 2533 1405 2556
rect 1430 2506 1433 2573
rect 1442 2513 1445 2643
rect 1450 2613 1453 2636
rect 1458 2586 1461 2726
rect 1466 2706 1469 2766
rect 1474 2723 1477 2826
rect 1482 2793 1485 2873
rect 1482 2733 1485 2746
rect 1490 2716 1493 2846
rect 1486 2713 1493 2716
rect 1466 2703 1473 2706
rect 1470 2646 1473 2703
rect 1486 2656 1489 2713
rect 1498 2663 1501 2986
rect 1510 2896 1513 2993
rect 1546 2983 1549 3040
rect 1570 2976 1573 3040
rect 1554 2973 1573 2976
rect 1586 2973 1589 3040
rect 1554 2953 1557 2973
rect 1626 2966 1629 3040
rect 1562 2963 1605 2966
rect 1522 2943 1557 2946
rect 1554 2926 1557 2943
rect 1562 2933 1565 2963
rect 1522 2923 1541 2926
rect 1554 2923 1565 2926
rect 1506 2893 1513 2896
rect 1506 2873 1509 2893
rect 1506 2733 1509 2776
rect 1546 2763 1549 2806
rect 1554 2746 1557 2816
rect 1562 2796 1565 2923
rect 1578 2886 1581 2936
rect 1602 2923 1605 2963
rect 1618 2963 1629 2966
rect 1642 2966 1645 3040
rect 1642 2963 1649 2966
rect 1618 2906 1621 2963
rect 1618 2903 1629 2906
rect 1578 2883 1613 2886
rect 1562 2793 1573 2796
rect 1570 2766 1573 2793
rect 1578 2773 1581 2816
rect 1586 2766 1589 2786
rect 1594 2776 1597 2806
rect 1610 2793 1613 2883
rect 1626 2843 1629 2903
rect 1646 2886 1649 2963
rect 1658 2923 1661 3040
rect 1674 2963 1677 3040
rect 1690 2983 1693 3040
rect 1706 2976 1709 3040
rect 1706 2973 1713 2976
rect 1642 2883 1649 2886
rect 1634 2776 1637 2816
rect 1642 2813 1645 2883
rect 1674 2856 1677 2936
rect 1658 2853 1677 2856
rect 1594 2773 1637 2776
rect 1570 2763 1605 2766
rect 1554 2743 1565 2746
rect 1602 2743 1605 2763
rect 1466 2643 1473 2646
rect 1482 2653 1489 2656
rect 1466 2593 1469 2643
rect 1482 2613 1485 2653
rect 1506 2643 1509 2726
rect 1554 2723 1557 2736
rect 1562 2703 1565 2743
rect 1578 2723 1605 2726
rect 1602 2706 1605 2723
rect 1598 2703 1605 2706
rect 1458 2583 1469 2586
rect 1466 2536 1469 2583
rect 1482 2553 1485 2606
rect 1506 2546 1509 2616
rect 1498 2543 1509 2546
rect 1466 2533 1493 2536
rect 1394 2476 1397 2506
rect 1426 2503 1433 2506
rect 1338 2463 1357 2466
rect 1370 2473 1377 2476
rect 1386 2473 1397 2476
rect 1338 2406 1341 2463
rect 1330 2403 1341 2406
rect 1270 2353 1277 2356
rect 1122 2216 1125 2233
rect 1138 2223 1141 2233
rect 1146 2216 1149 2226
rect 1122 2213 1149 2216
rect 1090 2203 1101 2206
rect 1090 2116 1093 2203
rect 1130 2133 1149 2136
rect 1090 2113 1101 2116
rect 1106 2113 1109 2126
rect 1026 2103 1061 2106
rect 994 2013 1005 2016
rect 962 1923 965 1936
rect 978 1933 989 1936
rect 938 1833 949 1836
rect 938 1786 941 1833
rect 946 1813 949 1826
rect 954 1803 957 1836
rect 938 1783 949 1786
rect 946 1726 949 1783
rect 962 1733 965 1746
rect 938 1723 949 1726
rect 914 1703 925 1706
rect 882 1623 885 1656
rect 906 1636 909 1696
rect 902 1633 909 1636
rect 890 1613 893 1626
rect 882 1593 885 1606
rect 890 1523 893 1586
rect 902 1566 905 1633
rect 922 1626 925 1703
rect 938 1676 941 1723
rect 914 1623 925 1626
rect 934 1673 941 1676
rect 934 1626 937 1673
rect 934 1623 941 1626
rect 914 1576 917 1623
rect 922 1603 933 1606
rect 914 1573 921 1576
rect 902 1563 909 1566
rect 906 1533 909 1563
rect 918 1526 921 1573
rect 914 1523 921 1526
rect 914 1506 917 1523
rect 906 1503 917 1506
rect 906 1426 909 1503
rect 906 1423 917 1426
rect 914 1406 917 1423
rect 930 1413 933 1516
rect 938 1406 941 1623
rect 946 1603 949 1666
rect 954 1523 957 1626
rect 962 1596 965 1716
rect 970 1606 973 1736
rect 978 1643 981 1926
rect 1002 1913 1005 2013
rect 1010 2043 1021 2046
rect 1010 1906 1013 2043
rect 1026 1983 1029 2103
rect 1098 2086 1101 2113
rect 1098 2083 1117 2086
rect 1074 2013 1077 2026
rect 1106 1993 1109 2016
rect 1114 2013 1117 2083
rect 1130 2076 1133 2133
rect 1146 2096 1149 2126
rect 1154 2123 1157 2233
rect 1146 2093 1173 2096
rect 1130 2073 1141 2076
rect 1138 2026 1141 2073
rect 1130 2023 1141 2026
rect 1018 1946 1021 1966
rect 1018 1943 1025 1946
rect 1002 1903 1013 1906
rect 994 1716 997 1726
rect 986 1713 997 1716
rect 994 1613 997 1636
rect 970 1603 981 1606
rect 962 1593 973 1596
rect 946 1413 949 1506
rect 962 1413 965 1586
rect 970 1556 973 1593
rect 978 1576 981 1603
rect 1002 1593 1005 1903
rect 1022 1896 1025 1943
rect 1018 1893 1025 1896
rect 1010 1813 1013 1836
rect 1018 1806 1021 1893
rect 1034 1816 1037 1956
rect 1058 1913 1061 1926
rect 1074 1826 1077 1976
rect 1082 1913 1085 1926
rect 1010 1803 1021 1806
rect 1026 1813 1037 1816
rect 1026 1796 1029 1813
rect 1042 1806 1045 1826
rect 1074 1823 1081 1826
rect 1018 1793 1029 1796
rect 1018 1723 1021 1793
rect 1034 1783 1037 1806
rect 1042 1803 1053 1806
rect 1050 1756 1053 1803
rect 1042 1753 1053 1756
rect 978 1573 989 1576
rect 970 1553 977 1556
rect 974 1476 977 1553
rect 970 1473 977 1476
rect 890 1373 893 1406
rect 906 1403 917 1406
rect 858 1363 877 1366
rect 842 1343 853 1346
rect 834 1333 845 1336
rect 794 1313 829 1316
rect 826 1226 829 1313
rect 770 1213 773 1226
rect 826 1223 837 1226
rect 834 1203 837 1223
rect 754 1113 757 1166
rect 714 1103 733 1106
rect 698 1053 709 1056
rect 690 1023 693 1036
rect 674 1013 701 1016
rect 706 1006 709 1053
rect 698 1003 709 1006
rect 674 913 677 936
rect 698 886 701 1003
rect 730 996 733 1103
rect 778 1006 781 1076
rect 810 1073 813 1126
rect 818 1123 821 1166
rect 842 1133 845 1333
rect 850 1196 853 1343
rect 858 1333 861 1363
rect 906 1356 909 1403
rect 906 1353 917 1356
rect 866 1333 901 1336
rect 858 1323 877 1326
rect 858 1306 861 1323
rect 858 1303 869 1306
rect 866 1236 869 1303
rect 858 1233 869 1236
rect 858 1213 861 1233
rect 882 1203 885 1333
rect 890 1323 901 1326
rect 906 1313 909 1326
rect 914 1296 917 1353
rect 922 1323 925 1406
rect 938 1403 949 1406
rect 906 1293 917 1296
rect 946 1296 949 1403
rect 970 1396 973 1473
rect 986 1456 989 1573
rect 978 1453 989 1456
rect 978 1406 981 1453
rect 994 1406 997 1436
rect 1002 1413 1005 1426
rect 978 1403 989 1406
rect 994 1403 1005 1406
rect 1010 1403 1013 1616
rect 1026 1613 1029 1736
rect 1034 1733 1037 1746
rect 1042 1723 1045 1753
rect 1066 1746 1069 1816
rect 1078 1776 1081 1823
rect 1098 1783 1101 1986
rect 1130 1883 1133 2023
rect 1162 2003 1165 2026
rect 1170 1963 1173 2093
rect 1178 1993 1181 2006
rect 1186 1986 1189 2316
rect 1202 2233 1205 2276
rect 1242 2206 1245 2226
rect 1234 2203 1245 2206
rect 1234 2136 1237 2203
rect 1258 2173 1261 2336
rect 1270 2286 1273 2353
rect 1282 2343 1309 2346
rect 1282 2313 1285 2343
rect 1270 2283 1277 2286
rect 1274 2233 1277 2283
rect 1290 2236 1293 2336
rect 1306 2313 1309 2343
rect 1322 2296 1325 2336
rect 1282 2233 1293 2236
rect 1314 2293 1325 2296
rect 1194 2113 1197 2136
rect 1202 2093 1205 2136
rect 1234 2133 1245 2136
rect 1226 2046 1229 2116
rect 1218 2043 1229 2046
rect 1194 2003 1197 2036
rect 1178 1983 1189 1986
rect 1146 1923 1149 1946
rect 1162 1926 1165 1936
rect 1178 1933 1181 1983
rect 1154 1923 1165 1926
rect 1218 1923 1221 2043
rect 1226 2013 1229 2036
rect 1242 2016 1245 2133
rect 1258 2123 1261 2136
rect 1234 2013 1245 2016
rect 1258 2013 1261 2026
rect 1226 1923 1229 1936
rect 1078 1773 1085 1776
rect 1066 1743 1073 1746
rect 1026 1533 1029 1556
rect 1034 1536 1037 1606
rect 1034 1533 1045 1536
rect 1026 1413 1029 1456
rect 1034 1426 1037 1526
rect 1050 1523 1053 1716
rect 1058 1693 1061 1736
rect 1070 1686 1073 1743
rect 1066 1683 1073 1686
rect 1066 1636 1069 1683
rect 1062 1633 1069 1636
rect 1062 1576 1065 1633
rect 1074 1603 1077 1626
rect 1062 1573 1069 1576
rect 1066 1553 1069 1573
rect 1074 1533 1077 1596
rect 1082 1573 1085 1773
rect 1098 1723 1101 1756
rect 1106 1733 1109 1746
rect 1114 1723 1117 1736
rect 1122 1706 1125 1736
rect 1114 1703 1125 1706
rect 1114 1646 1117 1703
rect 1114 1643 1125 1646
rect 1098 1613 1101 1636
rect 1122 1623 1125 1643
rect 1034 1423 1053 1426
rect 970 1393 981 1396
rect 978 1323 981 1393
rect 986 1323 989 1403
rect 1002 1333 1005 1403
rect 1034 1393 1037 1406
rect 1050 1333 1053 1423
rect 1074 1406 1077 1526
rect 1082 1413 1085 1426
rect 1074 1403 1085 1406
rect 1002 1303 1005 1326
rect 1066 1313 1069 1326
rect 946 1293 957 1296
rect 850 1193 885 1196
rect 858 1133 877 1136
rect 786 1013 789 1026
rect 778 1003 797 1006
rect 714 993 733 996
rect 714 923 717 993
rect 722 913 725 946
rect 730 913 733 936
rect 778 923 781 956
rect 850 946 853 1126
rect 882 1123 885 1193
rect 906 1136 909 1293
rect 930 1206 933 1286
rect 954 1226 957 1293
rect 1010 1226 1013 1246
rect 922 1203 933 1206
rect 946 1223 957 1226
rect 946 1203 949 1223
rect 986 1213 989 1226
rect 1010 1223 1021 1226
rect 922 1156 925 1203
rect 922 1153 929 1156
rect 906 1133 917 1136
rect 890 1073 893 1116
rect 914 1036 917 1133
rect 926 1096 929 1153
rect 938 1123 941 1196
rect 962 1193 973 1196
rect 1002 1183 1005 1216
rect 1018 1176 1021 1223
rect 1042 1203 1045 1216
rect 1058 1213 1069 1216
rect 1058 1206 1061 1213
rect 1050 1203 1061 1206
rect 1002 1133 1005 1176
rect 1010 1173 1021 1176
rect 962 1123 973 1126
rect 926 1093 933 1096
rect 930 1076 933 1093
rect 930 1073 957 1076
rect 914 1033 933 1036
rect 890 1013 893 1026
rect 930 983 933 1033
rect 954 1006 957 1073
rect 978 1066 981 1126
rect 1010 1106 1013 1173
rect 1034 1133 1037 1156
rect 1050 1126 1053 1203
rect 1074 1166 1077 1326
rect 1082 1303 1085 1403
rect 1090 1386 1093 1406
rect 1098 1403 1101 1606
rect 1114 1583 1117 1616
rect 1130 1613 1133 1876
rect 1154 1866 1157 1923
rect 1186 1913 1221 1916
rect 1146 1863 1157 1866
rect 1146 1813 1149 1863
rect 1186 1826 1189 1886
rect 1186 1823 1193 1826
rect 1138 1693 1141 1736
rect 1146 1613 1149 1636
rect 1122 1536 1125 1606
rect 1114 1533 1125 1536
rect 1146 1533 1149 1566
rect 1154 1533 1157 1556
rect 1090 1383 1097 1386
rect 1094 1296 1097 1383
rect 1090 1293 1097 1296
rect 1082 1203 1085 1246
rect 1090 1233 1093 1293
rect 1106 1226 1109 1416
rect 1114 1403 1117 1533
rect 1162 1526 1165 1776
rect 1178 1733 1181 1816
rect 1190 1756 1193 1823
rect 1186 1753 1193 1756
rect 1186 1733 1189 1753
rect 1202 1726 1205 1826
rect 1218 1813 1221 1913
rect 1234 1906 1237 2013
rect 1250 1933 1253 2006
rect 1230 1903 1237 1906
rect 1230 1836 1233 1903
rect 1230 1833 1237 1836
rect 1234 1813 1237 1833
rect 1242 1796 1245 1916
rect 1234 1793 1245 1796
rect 1210 1733 1213 1746
rect 1202 1723 1213 1726
rect 1186 1606 1189 1646
rect 1202 1613 1205 1626
rect 1186 1603 1197 1606
rect 1122 1413 1125 1426
rect 1138 1403 1141 1526
rect 1154 1523 1165 1526
rect 1154 1333 1157 1523
rect 1170 1513 1173 1526
rect 1194 1456 1197 1603
rect 1194 1453 1205 1456
rect 1170 1333 1173 1416
rect 1186 1403 1189 1436
rect 1202 1403 1205 1453
rect 1210 1386 1213 1723
rect 1218 1613 1221 1676
rect 1234 1636 1237 1793
rect 1234 1633 1245 1636
rect 1218 1526 1221 1606
rect 1242 1546 1245 1633
rect 1250 1556 1253 1926
rect 1258 1923 1261 1946
rect 1266 1906 1269 2216
rect 1282 2213 1285 2233
rect 1314 2226 1317 2293
rect 1314 2223 1325 2226
rect 1262 1903 1269 1906
rect 1262 1826 1265 1903
rect 1262 1823 1269 1826
rect 1258 1696 1261 1806
rect 1266 1716 1269 1823
rect 1274 1813 1277 2206
rect 1282 2203 1293 2206
rect 1282 2036 1285 2136
rect 1290 2123 1293 2176
rect 1298 2133 1301 2146
rect 1306 2133 1309 2206
rect 1314 2133 1317 2156
rect 1322 2116 1325 2223
rect 1314 2113 1325 2116
rect 1314 2056 1317 2113
rect 1314 2053 1325 2056
rect 1282 2033 1309 2036
rect 1282 2003 1285 2016
rect 1298 2013 1301 2026
rect 1282 1906 1285 1936
rect 1298 1933 1301 2006
rect 1306 2003 1309 2033
rect 1290 1923 1301 1926
rect 1306 1923 1309 1946
rect 1314 1923 1317 2016
rect 1322 1923 1325 2053
rect 1330 1906 1333 2403
rect 1370 2376 1373 2473
rect 1370 2373 1381 2376
rect 1378 2353 1381 2373
rect 1354 2343 1381 2346
rect 1338 2296 1341 2316
rect 1338 2293 1345 2296
rect 1342 1956 1345 2293
rect 1282 1903 1293 1906
rect 1274 1723 1277 1806
rect 1290 1796 1293 1903
rect 1322 1903 1333 1906
rect 1338 1953 1345 1956
rect 1322 1846 1325 1903
rect 1322 1843 1333 1846
rect 1306 1803 1309 1826
rect 1330 1823 1333 1843
rect 1282 1793 1293 1796
rect 1282 1773 1285 1793
rect 1266 1713 1277 1716
rect 1282 1713 1285 1726
rect 1258 1693 1265 1696
rect 1262 1636 1265 1693
rect 1258 1633 1265 1636
rect 1258 1603 1261 1633
rect 1274 1556 1277 1713
rect 1306 1666 1309 1786
rect 1330 1723 1333 1806
rect 1338 1706 1341 1953
rect 1346 1906 1349 1936
rect 1354 1926 1357 2343
rect 1362 2323 1365 2336
rect 1378 2333 1381 2343
rect 1386 2323 1389 2473
rect 1402 2456 1405 2496
rect 1426 2486 1429 2503
rect 1398 2453 1405 2456
rect 1410 2483 1429 2486
rect 1398 2376 1401 2453
rect 1410 2386 1413 2483
rect 1442 2423 1445 2436
rect 1426 2413 1445 2416
rect 1418 2403 1429 2406
rect 1450 2403 1453 2526
rect 1482 2523 1485 2533
rect 1466 2456 1469 2476
rect 1462 2453 1469 2456
rect 1410 2383 1421 2386
rect 1398 2373 1405 2376
rect 1402 2323 1405 2373
rect 1362 2313 1405 2316
rect 1418 2306 1421 2383
rect 1462 2356 1465 2453
rect 1442 2333 1445 2356
rect 1462 2353 1469 2356
rect 1410 2303 1421 2306
rect 1410 2263 1413 2303
rect 1466 2286 1469 2353
rect 1462 2283 1469 2286
rect 1378 2253 1421 2256
rect 1378 2213 1381 2253
rect 1418 2213 1421 2253
rect 1462 2206 1465 2283
rect 1474 2213 1477 2516
rect 1482 2316 1485 2466
rect 1490 2403 1493 2526
rect 1498 2496 1501 2543
rect 1522 2533 1525 2596
rect 1498 2493 1517 2496
rect 1498 2403 1501 2476
rect 1490 2323 1493 2346
rect 1506 2333 1509 2416
rect 1514 2406 1517 2493
rect 1522 2473 1525 2526
rect 1514 2403 1525 2406
rect 1522 2323 1525 2356
rect 1530 2316 1533 2666
rect 1598 2636 1601 2703
rect 1610 2663 1613 2716
rect 1598 2633 1605 2636
rect 1562 2593 1565 2616
rect 1570 2603 1573 2626
rect 1602 2613 1605 2633
rect 1634 2626 1637 2726
rect 1642 2713 1645 2736
rect 1658 2733 1661 2853
rect 1698 2836 1701 2966
rect 1710 2856 1713 2973
rect 1730 2963 1733 3040
rect 1746 2993 1749 3040
rect 1762 2986 1765 3040
rect 1722 2923 1725 2946
rect 1710 2853 1733 2856
rect 1674 2833 1701 2836
rect 1674 2746 1677 2833
rect 1682 2813 1693 2816
rect 1706 2803 1709 2816
rect 1730 2776 1733 2853
rect 1706 2773 1733 2776
rect 1674 2743 1693 2746
rect 1682 2713 1685 2726
rect 1690 2676 1693 2743
rect 1626 2623 1637 2626
rect 1682 2673 1693 2676
rect 1546 2556 1549 2586
rect 1626 2583 1629 2606
rect 1634 2573 1637 2606
rect 1650 2576 1653 2616
rect 1682 2576 1685 2673
rect 1698 2656 1701 2706
rect 1694 2653 1701 2656
rect 1694 2596 1697 2653
rect 1694 2593 1701 2596
rect 1650 2573 1661 2576
rect 1682 2573 1693 2576
rect 1538 2553 1549 2556
rect 1610 2563 1653 2566
rect 1538 2353 1541 2553
rect 1546 2393 1549 2546
rect 1610 2533 1613 2563
rect 1570 2523 1589 2526
rect 1626 2486 1629 2536
rect 1650 2523 1653 2563
rect 1658 2503 1661 2573
rect 1554 2386 1557 2486
rect 1618 2483 1629 2486
rect 1562 2413 1565 2436
rect 1578 2403 1581 2416
rect 1602 2403 1605 2426
rect 1562 2393 1597 2396
rect 1554 2383 1589 2386
rect 1546 2343 1565 2346
rect 1538 2323 1541 2336
rect 1546 2333 1549 2343
rect 1562 2326 1565 2343
rect 1570 2333 1573 2346
rect 1578 2333 1581 2356
rect 1562 2323 1573 2326
rect 1482 2313 1493 2316
rect 1394 2166 1397 2206
rect 1462 2203 1469 2206
rect 1482 2203 1485 2236
rect 1386 2163 1397 2166
rect 1386 2133 1389 2163
rect 1370 2106 1373 2126
rect 1370 2103 1389 2106
rect 1370 2013 1373 2036
rect 1386 2013 1389 2103
rect 1378 1976 1381 2006
rect 1402 2003 1405 2026
rect 1418 2013 1421 2126
rect 1466 2123 1469 2203
rect 1490 2103 1493 2313
rect 1514 2313 1533 2316
rect 1514 2246 1517 2313
rect 1570 2253 1573 2316
rect 1506 2243 1517 2246
rect 1506 2226 1509 2243
rect 1502 2223 1509 2226
rect 1502 2116 1505 2223
rect 1514 2123 1517 2186
rect 1554 2176 1557 2236
rect 1562 2183 1565 2216
rect 1586 2203 1589 2383
rect 1594 2343 1597 2393
rect 1618 2376 1621 2483
rect 1690 2476 1693 2573
rect 1686 2473 1693 2476
rect 1642 2413 1645 2426
rect 1618 2373 1661 2376
rect 1554 2173 1565 2176
rect 1502 2113 1509 2116
rect 1506 2096 1509 2113
rect 1514 2103 1517 2116
rect 1506 2093 1549 2096
rect 1434 2003 1437 2036
rect 1498 2023 1541 2026
rect 1474 2003 1485 2006
rect 1490 2003 1493 2016
rect 1498 2006 1501 2023
rect 1546 2006 1549 2093
rect 1498 2003 1509 2006
rect 1378 1973 1389 1976
rect 1386 1933 1389 1973
rect 1450 1963 1493 1966
rect 1354 1923 1381 1926
rect 1394 1923 1397 1936
rect 1346 1903 1357 1906
rect 1410 1903 1413 1936
rect 1450 1923 1453 1963
rect 1354 1776 1357 1903
rect 1370 1813 1373 1826
rect 1418 1813 1421 1826
rect 1298 1663 1309 1666
rect 1334 1703 1341 1706
rect 1350 1773 1357 1776
rect 1394 1776 1397 1806
rect 1466 1776 1469 1936
rect 1490 1923 1493 1963
rect 1506 1916 1509 2003
rect 1538 2003 1549 2006
rect 1538 1946 1541 2003
rect 1538 1943 1549 1946
rect 1546 1923 1549 1943
rect 1498 1913 1509 1916
rect 1482 1813 1485 1896
rect 1498 1856 1501 1913
rect 1494 1853 1501 1856
rect 1494 1806 1497 1853
rect 1394 1773 1469 1776
rect 1474 1803 1497 1806
rect 1282 1623 1285 1646
rect 1282 1576 1285 1606
rect 1298 1603 1301 1663
rect 1322 1576 1325 1616
rect 1282 1573 1325 1576
rect 1250 1553 1261 1556
rect 1274 1553 1285 1556
rect 1242 1543 1253 1546
rect 1218 1523 1225 1526
rect 1222 1466 1225 1523
rect 1218 1463 1225 1466
rect 1218 1433 1221 1463
rect 1202 1383 1213 1386
rect 1202 1326 1205 1383
rect 1218 1363 1221 1406
rect 1226 1336 1229 1446
rect 1234 1423 1237 1526
rect 1242 1523 1245 1536
rect 1250 1533 1253 1543
rect 1258 1536 1261 1553
rect 1258 1533 1265 1536
rect 1250 1503 1253 1526
rect 1262 1476 1265 1533
rect 1282 1486 1285 1553
rect 1314 1533 1317 1546
rect 1334 1516 1337 1703
rect 1350 1696 1353 1773
rect 1394 1763 1397 1773
rect 1386 1723 1389 1746
rect 1426 1733 1429 1773
rect 1474 1756 1477 1803
rect 1466 1753 1477 1756
rect 1346 1693 1353 1696
rect 1346 1533 1349 1693
rect 1378 1603 1381 1616
rect 1394 1613 1397 1646
rect 1258 1473 1265 1476
rect 1274 1483 1285 1486
rect 1330 1513 1337 1516
rect 1258 1456 1261 1473
rect 1250 1453 1261 1456
rect 1250 1376 1253 1453
rect 1266 1413 1269 1446
rect 1274 1413 1277 1483
rect 1282 1413 1293 1416
rect 1282 1393 1285 1413
rect 1298 1383 1301 1466
rect 1330 1446 1333 1513
rect 1346 1503 1349 1526
rect 1354 1453 1357 1526
rect 1370 1506 1373 1526
rect 1366 1503 1373 1506
rect 1306 1413 1309 1446
rect 1330 1443 1341 1446
rect 1250 1373 1293 1376
rect 1226 1333 1261 1336
rect 1122 1296 1125 1326
rect 1122 1293 1133 1296
rect 1130 1246 1133 1293
rect 1090 1223 1109 1226
rect 1122 1243 1133 1246
rect 1122 1223 1125 1243
rect 1162 1226 1165 1326
rect 1178 1313 1181 1326
rect 1202 1323 1213 1326
rect 1210 1226 1213 1323
rect 1234 1253 1237 1326
rect 1242 1323 1269 1326
rect 1066 1163 1077 1166
rect 1066 1146 1069 1163
rect 1018 1123 1053 1126
rect 1058 1143 1069 1146
rect 1058 1106 1061 1143
rect 1090 1133 1093 1223
rect 1010 1103 1029 1106
rect 970 1063 981 1066
rect 970 1013 973 1063
rect 1026 1036 1029 1103
rect 1050 1103 1061 1106
rect 1026 1033 1037 1036
rect 954 1003 965 1006
rect 802 943 829 946
rect 698 883 725 886
rect 642 793 645 806
rect 642 743 645 756
rect 378 673 397 676
rect 354 643 365 646
rect 282 593 293 596
rect 282 506 285 593
rect 306 533 309 586
rect 346 566 349 616
rect 362 583 365 643
rect 346 563 381 566
rect 282 503 293 506
rect 290 483 293 503
rect 298 373 325 376
rect 218 333 221 346
rect 274 206 277 336
rect 298 333 301 373
rect 282 316 285 326
rect 306 323 309 366
rect 314 316 317 336
rect 322 333 325 373
rect 330 316 333 416
rect 354 413 357 526
rect 354 383 357 406
rect 370 363 373 416
rect 282 313 317 316
rect 322 313 333 316
rect 322 296 325 313
rect 314 293 325 296
rect 314 236 317 293
rect 314 233 325 236
rect 274 203 285 206
rect 258 73 261 196
rect 282 146 285 203
rect 322 196 325 233
rect 274 143 285 146
rect 314 193 325 196
rect 274 123 277 143
rect 314 136 317 193
rect 314 133 325 136
rect 322 103 325 133
rect 330 123 333 136
rect 2 3 85 6
rect 338 0 341 336
rect 346 266 349 336
rect 346 263 365 266
rect 362 206 365 263
rect 378 226 381 563
rect 386 523 389 536
rect 394 533 397 673
rect 410 576 413 616
rect 442 613 445 646
rect 458 643 461 726
rect 466 703 469 726
rect 482 723 493 726
rect 410 573 453 576
rect 450 536 453 573
rect 418 516 421 536
rect 450 533 461 536
rect 410 513 421 516
rect 410 446 413 513
rect 434 453 437 526
rect 458 523 461 533
rect 482 506 485 723
rect 506 613 509 726
rect 562 706 565 726
rect 562 703 573 706
rect 546 676 549 696
rect 538 673 549 676
rect 538 626 541 673
rect 570 636 573 703
rect 562 633 573 636
rect 538 623 549 626
rect 474 503 485 506
rect 474 456 477 503
rect 474 453 485 456
rect 410 443 421 446
rect 418 423 421 443
rect 482 433 485 453
rect 498 423 501 606
rect 546 603 549 623
rect 562 613 565 633
rect 610 613 613 646
rect 618 616 621 736
rect 690 733 693 816
rect 722 813 725 883
rect 738 793 741 806
rect 730 743 741 746
rect 634 693 637 716
rect 706 706 709 726
rect 690 703 709 706
rect 634 623 653 626
rect 618 613 653 616
rect 554 533 557 546
rect 570 533 573 586
rect 482 413 493 416
rect 426 343 429 406
rect 410 333 429 336
rect 402 306 405 326
rect 394 303 405 306
rect 394 256 397 303
rect 394 253 405 256
rect 378 223 385 226
rect 354 203 365 206
rect 354 126 357 203
rect 370 133 373 216
rect 382 126 385 223
rect 394 133 397 236
rect 402 216 405 253
rect 410 223 413 296
rect 426 286 429 333
rect 442 293 445 346
rect 458 323 461 336
rect 474 316 477 406
rect 490 396 493 413
rect 490 393 501 396
rect 498 333 501 393
rect 506 383 509 406
rect 506 323 509 346
rect 522 333 525 526
rect 602 523 605 546
rect 634 516 637 606
rect 650 523 653 613
rect 690 546 693 703
rect 690 543 709 546
rect 658 516 661 536
rect 706 523 709 543
rect 714 516 717 736
rect 738 616 741 743
rect 738 613 757 616
rect 762 613 765 746
rect 786 733 789 816
rect 818 813 821 926
rect 826 903 829 943
rect 842 943 853 946
rect 866 943 869 956
rect 834 913 837 936
rect 842 916 845 943
rect 850 933 893 936
rect 842 913 885 916
rect 874 826 877 906
rect 890 903 893 933
rect 874 823 885 826
rect 834 793 837 806
rect 794 743 813 746
rect 810 733 813 743
rect 794 723 813 726
rect 842 716 845 736
rect 834 713 845 716
rect 834 606 837 713
rect 858 656 861 726
rect 874 723 877 816
rect 882 776 885 823
rect 882 773 893 776
rect 890 736 893 773
rect 886 733 893 736
rect 886 676 889 733
rect 898 676 901 956
rect 938 923 941 936
rect 906 896 909 916
rect 906 893 917 896
rect 914 836 917 893
rect 954 876 957 926
rect 962 913 965 1003
rect 1010 953 1013 1016
rect 1018 1003 1021 1026
rect 1034 986 1037 1033
rect 1026 983 1037 986
rect 1002 903 1005 926
rect 954 873 961 876
rect 906 833 917 836
rect 906 693 909 833
rect 946 816 949 866
rect 958 826 961 873
rect 1018 863 1021 936
rect 1026 933 1029 983
rect 1050 966 1053 1103
rect 1042 963 1053 966
rect 1042 946 1045 963
rect 1066 956 1069 1126
rect 1082 963 1085 1016
rect 1038 943 1045 946
rect 1050 953 1069 956
rect 1038 866 1041 943
rect 1038 863 1045 866
rect 914 753 917 816
rect 922 813 949 816
rect 954 823 961 826
rect 938 793 941 806
rect 954 786 957 823
rect 922 783 957 786
rect 886 673 893 676
rect 898 673 905 676
rect 858 653 885 656
rect 786 593 789 606
rect 794 583 797 606
rect 834 603 845 606
rect 842 586 845 603
rect 858 586 861 606
rect 882 593 885 653
rect 890 586 893 673
rect 802 583 861 586
rect 770 533 773 576
rect 634 513 661 516
rect 698 513 717 516
rect 714 466 717 513
rect 714 463 725 466
rect 474 313 525 316
rect 538 313 541 416
rect 650 413 653 456
rect 546 363 549 406
rect 546 333 581 336
rect 426 283 445 286
rect 402 213 421 216
rect 418 146 421 213
rect 418 143 429 146
rect 354 123 365 126
rect 362 83 365 123
rect 378 123 385 126
rect 426 123 429 143
rect 378 73 381 123
rect 442 113 445 283
rect 490 203 493 296
rect 514 223 517 236
rect 498 213 517 216
rect 490 116 493 136
rect 506 123 509 213
rect 522 203 525 313
rect 546 206 549 316
rect 562 216 565 326
rect 578 313 581 333
rect 562 213 589 216
rect 546 203 573 206
rect 546 133 549 186
rect 554 133 557 146
rect 490 113 525 116
rect 474 86 477 106
rect 570 93 573 203
rect 586 103 589 206
rect 602 133 605 226
rect 618 203 621 406
rect 682 376 685 426
rect 722 413 725 463
rect 698 393 701 406
rect 778 383 781 416
rect 802 393 805 583
rect 818 563 861 566
rect 818 523 821 563
rect 858 533 861 563
rect 850 413 853 526
rect 866 456 869 546
rect 874 523 877 586
rect 886 583 893 586
rect 886 516 889 583
rect 902 576 905 673
rect 922 656 925 783
rect 962 733 965 806
rect 978 766 981 806
rect 1026 803 1029 816
rect 1042 806 1045 863
rect 1050 826 1053 953
rect 1058 843 1061 926
rect 1074 923 1077 936
rect 1098 923 1101 1006
rect 1114 916 1117 1216
rect 1130 1203 1133 1226
rect 1162 1223 1181 1226
rect 1210 1223 1245 1226
rect 1162 1196 1165 1216
rect 1154 1193 1165 1196
rect 1154 1146 1157 1193
rect 1154 1143 1165 1146
rect 1162 1126 1165 1143
rect 1178 1133 1181 1223
rect 1186 1193 1189 1216
rect 1210 1213 1237 1216
rect 1130 1083 1133 1116
rect 1138 966 1141 1126
rect 1162 1123 1197 1126
rect 1194 1086 1197 1123
rect 1178 1083 1197 1086
rect 1202 1083 1205 1206
rect 1210 1203 1213 1213
rect 1242 1206 1245 1223
rect 1226 1193 1229 1206
rect 1234 1203 1245 1206
rect 1250 1203 1253 1323
rect 1266 1313 1269 1323
rect 1290 1316 1293 1373
rect 1338 1346 1341 1443
rect 1366 1426 1369 1503
rect 1378 1463 1381 1536
rect 1386 1533 1389 1586
rect 1386 1503 1389 1526
rect 1418 1426 1421 1626
rect 1450 1613 1453 1726
rect 1466 1686 1469 1753
rect 1506 1723 1509 1846
rect 1554 1816 1557 2156
rect 1562 2116 1565 2173
rect 1562 2113 1569 2116
rect 1566 2046 1569 2113
rect 1578 2103 1581 2116
rect 1566 2043 1573 2046
rect 1562 1953 1565 2016
rect 1570 1993 1573 2043
rect 1602 2013 1605 2336
rect 1634 2333 1637 2346
rect 1658 2333 1661 2373
rect 1686 2356 1689 2473
rect 1698 2413 1701 2593
rect 1706 2523 1709 2773
rect 1738 2703 1741 2986
rect 1750 2983 1765 2986
rect 1750 2836 1753 2983
rect 1778 2976 1781 3040
rect 1802 2986 1805 3040
rect 1802 2983 1813 2986
rect 1762 2973 1781 2976
rect 1786 2973 1805 2976
rect 1762 2923 1765 2973
rect 1770 2933 1773 2946
rect 1778 2856 1781 2966
rect 1786 2943 1789 2973
rect 1802 2943 1805 2973
rect 1810 2936 1813 2983
rect 1746 2833 1753 2836
rect 1770 2853 1781 2856
rect 1794 2933 1813 2936
rect 1746 2723 1749 2833
rect 1754 2793 1757 2816
rect 1762 2733 1765 2746
rect 1714 2613 1717 2626
rect 1730 2613 1733 2686
rect 1754 2656 1757 2726
rect 1770 2716 1773 2853
rect 1738 2653 1757 2656
rect 1766 2713 1773 2716
rect 1706 2406 1709 2436
rect 1698 2403 1709 2406
rect 1714 2406 1717 2556
rect 1722 2513 1725 2606
rect 1730 2416 1733 2526
rect 1738 2503 1741 2653
rect 1746 2603 1749 2646
rect 1754 2613 1757 2626
rect 1766 2576 1769 2713
rect 1778 2586 1781 2846
rect 1786 2733 1789 2796
rect 1786 2683 1789 2716
rect 1778 2583 1785 2586
rect 1766 2573 1773 2576
rect 1770 2553 1773 2573
rect 1754 2533 1757 2546
rect 1782 2496 1785 2583
rect 1778 2493 1785 2496
rect 1730 2413 1757 2416
rect 1714 2403 1741 2406
rect 1698 2356 1701 2403
rect 1706 2373 1709 2396
rect 1686 2353 1693 2356
rect 1698 2353 1705 2356
rect 1626 2323 1645 2326
rect 1682 2323 1685 2336
rect 1690 2316 1693 2353
rect 1682 2313 1693 2316
rect 1682 2276 1685 2313
rect 1702 2306 1705 2353
rect 1738 2323 1741 2403
rect 1754 2333 1757 2346
rect 1770 2343 1773 2406
rect 1778 2363 1781 2493
rect 1786 2403 1789 2416
rect 1786 2323 1789 2346
rect 1674 2273 1685 2276
rect 1698 2303 1705 2306
rect 1618 2003 1621 2266
rect 1626 2233 1653 2236
rect 1626 2203 1629 2233
rect 1634 2223 1645 2226
rect 1626 2133 1629 2146
rect 1634 2123 1637 2216
rect 1650 2203 1653 2233
rect 1626 2013 1629 2036
rect 1626 1993 1629 2006
rect 1642 2003 1645 2106
rect 1650 2093 1653 2116
rect 1674 2036 1677 2273
rect 1698 2236 1701 2303
rect 1690 2233 1701 2236
rect 1690 2146 1693 2233
rect 1706 2156 1709 2226
rect 1746 2223 1757 2226
rect 1714 2203 1717 2216
rect 1706 2153 1713 2156
rect 1690 2143 1701 2146
rect 1698 2123 1701 2143
rect 1674 2033 1685 2036
rect 1666 1983 1669 2016
rect 1682 2006 1685 2033
rect 1698 2013 1701 2086
rect 1710 2026 1713 2153
rect 1722 2113 1725 2216
rect 1730 2136 1733 2216
rect 1730 2133 1757 2136
rect 1786 2133 1789 2146
rect 1730 2046 1733 2126
rect 1738 2063 1741 2106
rect 1746 2093 1749 2116
rect 1706 2023 1713 2026
rect 1722 2043 1733 2046
rect 1682 2003 1701 2006
rect 1602 1963 1645 1966
rect 1578 1933 1581 1946
rect 1602 1933 1605 1963
rect 1618 1933 1621 1946
rect 1554 1813 1561 1816
rect 1522 1726 1525 1806
rect 1466 1683 1477 1686
rect 1458 1603 1461 1626
rect 1474 1586 1477 1683
rect 1514 1676 1517 1726
rect 1522 1723 1533 1726
rect 1506 1673 1517 1676
rect 1474 1583 1481 1586
rect 1466 1556 1469 1576
rect 1450 1553 1469 1556
rect 1450 1446 1453 1553
rect 1478 1536 1481 1583
rect 1474 1533 1481 1536
rect 1450 1443 1469 1446
rect 1362 1423 1369 1426
rect 1362 1403 1365 1423
rect 1370 1363 1373 1416
rect 1378 1346 1381 1426
rect 1386 1403 1389 1426
rect 1402 1423 1437 1426
rect 1402 1356 1405 1423
rect 1402 1353 1413 1356
rect 1338 1343 1381 1346
rect 1338 1333 1341 1343
rect 1282 1313 1293 1316
rect 1282 1246 1285 1313
rect 1282 1243 1293 1246
rect 1290 1223 1293 1243
rect 1210 1123 1213 1136
rect 1234 1116 1237 1203
rect 1258 1173 1261 1216
rect 1274 1203 1277 1216
rect 1298 1196 1301 1326
rect 1322 1323 1349 1326
rect 1362 1323 1365 1336
rect 1410 1333 1413 1353
rect 1418 1346 1421 1416
rect 1426 1403 1437 1406
rect 1458 1386 1461 1406
rect 1418 1343 1429 1346
rect 1370 1313 1373 1326
rect 1418 1283 1421 1336
rect 1314 1246 1317 1266
rect 1290 1193 1301 1196
rect 1310 1243 1317 1246
rect 1310 1186 1313 1243
rect 1310 1183 1317 1186
rect 1250 1143 1261 1146
rect 1314 1133 1317 1183
rect 1218 1113 1237 1116
rect 1242 1113 1245 1126
rect 1258 1123 1269 1126
rect 1154 1003 1157 1016
rect 1138 963 1145 966
rect 1098 913 1117 916
rect 1050 823 1061 826
rect 1042 803 1049 806
rect 978 763 989 766
rect 970 723 973 746
rect 922 653 929 656
rect 926 576 929 653
rect 882 513 889 516
rect 898 573 905 576
rect 922 573 929 576
rect 866 453 873 456
rect 870 376 873 453
rect 682 373 709 376
rect 658 326 661 336
rect 634 323 661 326
rect 690 323 693 346
rect 706 333 709 373
rect 754 333 757 356
rect 626 143 629 316
rect 634 306 637 323
rect 634 303 645 306
rect 642 246 645 303
rect 634 243 645 246
rect 634 223 637 243
rect 658 196 661 323
rect 674 313 709 316
rect 674 223 693 226
rect 674 213 677 223
rect 682 196 685 216
rect 690 203 693 223
rect 658 193 685 196
rect 746 196 749 216
rect 746 193 757 196
rect 618 113 621 136
rect 650 126 653 146
rect 642 123 653 126
rect 466 83 477 86
rect 466 16 469 83
rect 466 13 477 16
rect 474 0 477 13
rect 490 0 493 86
rect 626 83 629 106
rect 506 0 509 76
rect 642 66 645 123
rect 658 73 661 186
rect 666 103 669 116
rect 674 93 677 126
rect 698 106 701 136
rect 738 123 741 136
rect 754 133 757 193
rect 762 123 765 376
rect 866 373 873 376
rect 778 333 781 346
rect 786 323 789 336
rect 778 293 781 316
rect 778 183 781 196
rect 722 113 757 116
rect 682 103 701 106
rect 770 73 773 136
rect 810 133 813 336
rect 842 333 845 356
rect 834 143 837 156
rect 826 123 829 136
rect 842 123 845 316
rect 866 223 869 373
rect 882 356 885 513
rect 890 373 893 416
rect 898 366 901 573
rect 922 536 925 573
rect 914 533 925 536
rect 914 376 917 533
rect 938 446 941 696
rect 986 686 989 763
rect 1010 733 1013 746
rect 970 683 989 686
rect 946 626 949 646
rect 946 623 953 626
rect 950 566 953 623
rect 970 586 973 683
rect 946 563 953 566
rect 962 583 973 586
rect 946 523 949 563
rect 962 533 965 583
rect 938 443 949 446
rect 946 396 949 443
rect 962 413 965 466
rect 986 413 989 526
rect 1002 426 1005 726
rect 1018 613 1021 736
rect 1034 643 1037 746
rect 1046 686 1049 803
rect 1042 683 1049 686
rect 1042 543 1045 683
rect 1058 566 1061 823
rect 1082 723 1085 806
rect 1050 563 1061 566
rect 1026 523 1045 526
rect 1002 423 1013 426
rect 994 396 997 416
rect 938 393 949 396
rect 990 393 997 396
rect 914 373 925 376
rect 878 353 885 356
rect 890 363 901 366
rect 878 286 881 353
rect 890 296 893 363
rect 890 293 901 296
rect 878 283 885 286
rect 882 216 885 283
rect 866 213 885 216
rect 858 133 861 146
rect 866 106 869 213
rect 898 206 901 293
rect 922 253 925 373
rect 938 346 941 393
rect 938 343 949 346
rect 946 286 949 343
rect 970 323 973 346
rect 990 336 993 393
rect 1010 366 1013 423
rect 1026 413 1029 523
rect 1050 516 1053 563
rect 1042 513 1053 516
rect 1042 406 1045 513
rect 1058 463 1061 536
rect 1066 526 1069 546
rect 1074 543 1077 646
rect 1066 523 1077 526
rect 1090 523 1093 736
rect 1098 723 1101 913
rect 1142 886 1145 963
rect 1138 883 1145 886
rect 1122 803 1133 806
rect 1138 753 1141 883
rect 1154 746 1157 926
rect 1178 856 1181 1083
rect 1202 1056 1205 1076
rect 1194 1053 1205 1056
rect 1194 986 1197 1053
rect 1218 1046 1221 1113
rect 1210 1043 1221 1046
rect 1194 983 1205 986
rect 1202 916 1205 983
rect 1210 933 1213 1043
rect 1218 1023 1245 1026
rect 1218 946 1221 1016
rect 1242 1013 1245 1023
rect 1258 1013 1261 1123
rect 1306 1093 1309 1126
rect 1330 1106 1333 1206
rect 1378 1193 1381 1216
rect 1402 1213 1413 1216
rect 1418 1206 1421 1226
rect 1410 1203 1421 1206
rect 1322 1103 1333 1106
rect 1226 993 1229 1006
rect 1234 1003 1245 1006
rect 1218 943 1237 946
rect 1210 923 1221 926
rect 1202 913 1221 916
rect 1218 856 1221 913
rect 1178 853 1197 856
rect 1218 853 1229 856
rect 1194 836 1197 853
rect 1194 833 1221 836
rect 1170 823 1189 826
rect 1186 816 1189 823
rect 1146 743 1157 746
rect 1106 733 1117 736
rect 1146 726 1149 743
rect 1138 723 1149 726
rect 1138 636 1141 723
rect 1154 706 1157 736
rect 1170 723 1173 816
rect 1178 803 1181 816
rect 1186 813 1197 816
rect 1202 733 1205 806
rect 1210 783 1213 806
rect 1186 716 1189 726
rect 1218 723 1221 833
rect 1226 813 1229 853
rect 1234 803 1237 943
rect 1266 923 1269 986
rect 1282 976 1285 1006
rect 1306 993 1309 1016
rect 1322 996 1325 1103
rect 1354 1016 1357 1136
rect 1410 1123 1413 1203
rect 1426 1146 1429 1343
rect 1442 1333 1445 1386
rect 1454 1383 1461 1386
rect 1454 1326 1457 1383
rect 1434 1203 1437 1326
rect 1450 1323 1457 1326
rect 1442 1173 1445 1216
rect 1426 1143 1433 1146
rect 1354 1013 1381 1016
rect 1322 993 1333 996
rect 1322 976 1325 993
rect 1282 973 1325 976
rect 1394 973 1397 1016
rect 1402 976 1405 1116
rect 1418 1106 1421 1136
rect 1414 1103 1421 1106
rect 1414 1036 1417 1103
rect 1430 1096 1433 1143
rect 1442 1113 1445 1126
rect 1410 1033 1417 1036
rect 1426 1093 1433 1096
rect 1410 1013 1413 1033
rect 1426 1013 1429 1093
rect 1410 983 1413 1006
rect 1426 993 1429 1006
rect 1402 973 1429 976
rect 1282 846 1285 973
rect 1322 933 1325 973
rect 1370 923 1373 956
rect 1402 886 1405 906
rect 1242 843 1285 846
rect 1242 786 1245 843
rect 1290 803 1293 816
rect 1242 783 1253 786
rect 1234 756 1237 776
rect 1230 753 1237 756
rect 1162 713 1189 716
rect 1230 706 1233 753
rect 1154 703 1165 706
rect 1230 703 1237 706
rect 1106 633 1141 636
rect 1106 586 1109 633
rect 1162 603 1165 703
rect 1106 583 1117 586
rect 1074 456 1077 523
rect 1098 506 1101 536
rect 1058 453 1077 456
rect 1090 503 1101 506
rect 986 333 993 336
rect 1002 363 1013 366
rect 1034 403 1045 406
rect 930 283 949 286
rect 882 203 901 206
rect 882 186 885 203
rect 858 103 869 106
rect 878 183 885 186
rect 642 63 653 66
rect 650 0 653 63
rect 858 16 861 103
rect 878 96 881 183
rect 930 156 933 283
rect 986 276 989 333
rect 978 273 989 276
rect 890 133 893 156
rect 922 153 933 156
rect 890 103 893 116
rect 922 106 925 153
rect 954 133 957 256
rect 978 216 981 273
rect 978 213 989 216
rect 978 123 981 196
rect 986 186 989 213
rect 994 193 997 206
rect 986 183 993 186
rect 922 103 933 106
rect 878 93 885 96
rect 858 13 869 16
rect 866 0 869 13
rect 882 0 885 93
rect 930 0 933 103
rect 978 76 981 116
rect 970 73 981 76
rect 990 76 993 183
rect 1002 86 1005 363
rect 1010 333 1013 346
rect 1034 326 1037 403
rect 1050 356 1053 406
rect 1058 366 1061 453
rect 1090 436 1093 503
rect 1114 436 1117 583
rect 1090 433 1101 436
rect 1082 403 1085 416
rect 1098 393 1101 433
rect 1110 433 1117 436
rect 1110 376 1113 433
rect 1122 423 1149 426
rect 1106 373 1113 376
rect 1058 363 1069 366
rect 1050 353 1061 356
rect 1018 113 1021 326
rect 1030 323 1037 326
rect 1058 323 1061 353
rect 1066 323 1069 363
rect 1030 226 1033 323
rect 1030 223 1037 226
rect 1034 203 1037 223
rect 1042 213 1045 316
rect 1074 313 1077 336
rect 1106 246 1109 373
rect 1130 343 1133 416
rect 1146 413 1149 423
rect 1138 396 1141 406
rect 1146 403 1157 406
rect 1178 396 1181 536
rect 1186 523 1189 626
rect 1202 563 1205 636
rect 1234 623 1237 703
rect 1250 686 1253 783
rect 1298 746 1301 836
rect 1322 813 1325 856
rect 1378 803 1381 886
rect 1394 883 1405 886
rect 1394 826 1397 883
rect 1394 823 1405 826
rect 1394 773 1397 806
rect 1402 756 1405 823
rect 1410 803 1413 926
rect 1290 743 1301 746
rect 1398 753 1405 756
rect 1250 683 1261 686
rect 1202 426 1205 536
rect 1250 533 1253 586
rect 1258 576 1261 683
rect 1258 573 1269 576
rect 1266 533 1269 573
rect 1290 546 1293 743
rect 1298 723 1301 736
rect 1330 713 1333 726
rect 1378 713 1381 726
rect 1386 693 1389 726
rect 1398 656 1401 753
rect 1410 733 1413 746
rect 1418 726 1421 966
rect 1410 723 1421 726
rect 1398 653 1405 656
rect 1306 603 1309 616
rect 1338 586 1341 616
rect 1394 613 1397 636
rect 1330 583 1341 586
rect 1290 543 1301 546
rect 1250 486 1253 526
rect 1298 486 1301 543
rect 1314 523 1317 546
rect 1250 483 1301 486
rect 1330 466 1333 583
rect 1338 523 1349 526
rect 1274 463 1333 466
rect 1202 423 1221 426
rect 1194 403 1197 416
rect 1202 413 1213 416
rect 1138 393 1181 396
rect 1202 383 1205 406
rect 1106 243 1117 246
rect 1106 213 1109 226
rect 1066 193 1069 206
rect 1050 153 1069 156
rect 1050 133 1053 153
rect 1066 133 1069 153
rect 1002 83 1013 86
rect 990 73 997 76
rect 970 16 973 73
rect 970 13 981 16
rect 978 0 981 13
rect 994 0 997 73
rect 1010 0 1013 83
rect 1034 0 1037 126
rect 1106 123 1109 146
rect 1114 53 1117 243
rect 1130 223 1133 336
rect 1186 333 1189 356
rect 1210 333 1213 413
rect 1194 316 1197 326
rect 1170 313 1197 316
rect 1178 213 1181 246
rect 1210 203 1213 226
rect 1154 133 1157 146
rect 1186 143 1189 156
rect 1146 66 1149 126
rect 1218 123 1221 423
rect 1226 393 1229 416
rect 1266 396 1269 416
rect 1274 403 1277 463
rect 1258 393 1269 396
rect 1258 346 1261 393
rect 1258 343 1269 346
rect 1266 323 1269 343
rect 1274 323 1277 346
rect 1282 316 1285 416
rect 1330 413 1333 436
rect 1354 413 1357 566
rect 1394 503 1397 526
rect 1402 486 1405 653
rect 1410 523 1413 723
rect 1418 703 1421 716
rect 1394 483 1405 486
rect 1394 406 1397 483
rect 1410 413 1413 426
rect 1290 343 1293 406
rect 1330 386 1333 406
rect 1394 403 1405 406
rect 1418 403 1421 646
rect 1426 526 1429 973
rect 1450 946 1453 1323
rect 1466 1296 1469 1443
rect 1474 1323 1477 1533
rect 1490 1426 1493 1626
rect 1506 1513 1509 1673
rect 1530 1666 1533 1723
rect 1522 1663 1533 1666
rect 1522 1603 1525 1663
rect 1546 1613 1549 1806
rect 1558 1716 1561 1813
rect 1570 1736 1573 1816
rect 1594 1803 1597 1926
rect 1642 1923 1645 1963
rect 1634 1803 1637 1816
rect 1666 1793 1669 1936
rect 1698 1923 1701 2003
rect 1706 1993 1709 2023
rect 1722 2013 1725 2043
rect 1730 2023 1733 2036
rect 1786 2033 1789 2116
rect 1794 1996 1797 2933
rect 1802 2906 1805 2926
rect 1802 2903 1813 2906
rect 1810 2846 1813 2903
rect 1802 2843 1813 2846
rect 1834 2843 1837 3040
rect 1954 3037 1973 3040
rect 1874 2963 1917 2966
rect 1874 2933 1877 2963
rect 1802 2733 1805 2843
rect 1818 2803 1821 2816
rect 1850 2696 1853 2736
rect 1842 2693 1853 2696
rect 1810 2613 1813 2686
rect 1826 2613 1829 2636
rect 1802 2583 1805 2606
rect 1802 2456 1805 2526
rect 1818 2503 1821 2606
rect 1802 2453 1813 2456
rect 1802 2423 1805 2436
rect 1810 2403 1813 2453
rect 1826 2386 1829 2586
rect 1842 2566 1845 2693
rect 1858 2603 1861 2926
rect 1890 2923 1893 2936
rect 1914 2923 1917 2963
rect 1954 2926 1957 3037
rect 2050 3026 2053 3040
rect 2042 3023 2053 3026
rect 2042 2976 2045 3023
rect 2042 2973 2053 2976
rect 1954 2923 1973 2926
rect 1986 2923 1989 2936
rect 2050 2926 2053 2973
rect 2066 2936 2069 3040
rect 2082 3026 2085 3040
rect 2082 3023 2093 3026
rect 2074 2943 2077 2956
rect 2066 2933 2077 2936
rect 2018 2913 2021 2926
rect 2050 2923 2069 2926
rect 1866 2776 1869 2816
rect 1914 2813 1917 2826
rect 1930 2803 1933 2816
rect 1866 2773 1901 2776
rect 1898 2733 1901 2773
rect 1874 2713 1877 2726
rect 1882 2723 1901 2726
rect 1882 2703 1885 2723
rect 1898 2683 1901 2716
rect 1906 2613 1909 2636
rect 1914 2613 1917 2626
rect 1938 2616 1941 2686
rect 1946 2666 1949 2776
rect 1978 2746 1981 2816
rect 2026 2773 2029 2816
rect 2050 2803 2053 2916
rect 2074 2886 2077 2933
rect 2066 2883 2077 2886
rect 2066 2826 2069 2883
rect 2090 2876 2093 3023
rect 2062 2823 2069 2826
rect 2082 2873 2093 2876
rect 2050 2783 2053 2796
rect 2062 2776 2065 2823
rect 2062 2773 2069 2776
rect 2074 2773 2077 2816
rect 2066 2756 2069 2773
rect 2066 2753 2073 2756
rect 1978 2743 1989 2746
rect 1986 2733 1989 2743
rect 2058 2733 2061 2746
rect 1986 2683 1989 2716
rect 1946 2663 1957 2666
rect 1930 2613 1941 2616
rect 1946 2613 1949 2656
rect 1906 2583 1909 2606
rect 1834 2563 1845 2566
rect 1922 2563 1925 2606
rect 1938 2593 1941 2606
rect 1954 2603 1957 2663
rect 2018 2633 2029 2636
rect 2042 2633 2045 2716
rect 2058 2686 2061 2726
rect 2054 2683 2061 2686
rect 2018 2623 2029 2626
rect 2018 2613 2021 2623
rect 2054 2616 2057 2683
rect 2070 2676 2073 2753
rect 2066 2673 2073 2676
rect 2066 2626 2069 2673
rect 2066 2623 2073 2626
rect 2050 2613 2057 2616
rect 1834 2513 1837 2563
rect 1858 2476 1861 2546
rect 1842 2473 1861 2476
rect 1906 2473 1909 2526
rect 1938 2523 1941 2566
rect 2018 2563 2021 2606
rect 1970 2506 1973 2526
rect 1962 2503 1973 2506
rect 1842 2403 1845 2473
rect 1962 2446 1965 2503
rect 1986 2486 1989 2536
rect 1986 2483 2005 2486
rect 1962 2443 1973 2446
rect 1826 2383 1845 2386
rect 1834 2323 1837 2366
rect 1842 2333 1845 2383
rect 1866 2236 1869 2436
rect 1874 2303 1877 2326
rect 1882 2323 1885 2416
rect 1890 2336 1893 2416
rect 1922 2403 1925 2416
rect 1954 2413 1957 2426
rect 1954 2383 1957 2406
rect 1970 2383 1973 2443
rect 1954 2343 1957 2366
rect 1890 2333 1901 2336
rect 1898 2283 1901 2316
rect 1970 2303 1973 2326
rect 1818 2203 1821 2236
rect 1802 2006 1805 2106
rect 1826 2063 1829 2236
rect 1862 2233 1869 2236
rect 1842 2126 1845 2226
rect 1850 2193 1853 2206
rect 1862 2176 1865 2233
rect 1862 2173 1869 2176
rect 1866 2153 1869 2173
rect 1842 2123 1861 2126
rect 1858 2113 1861 2123
rect 1866 2116 1869 2136
rect 1874 2133 1877 2146
rect 1914 2116 1917 2216
rect 1866 2113 1877 2116
rect 1834 2023 1837 2046
rect 1802 2003 1821 2006
rect 1794 1993 1805 1996
rect 1570 1733 1581 1736
rect 1650 1733 1669 1736
rect 1642 1723 1653 1726
rect 1658 1716 1661 1726
rect 1558 1713 1565 1716
rect 1634 1713 1661 1716
rect 1562 1636 1565 1713
rect 1558 1633 1565 1636
rect 1594 1633 1637 1636
rect 1546 1596 1549 1606
rect 1538 1593 1549 1596
rect 1538 1533 1541 1593
rect 1558 1586 1561 1633
rect 1554 1583 1561 1586
rect 1482 1423 1501 1426
rect 1482 1396 1485 1423
rect 1482 1393 1493 1396
rect 1482 1323 1485 1346
rect 1490 1313 1493 1393
rect 1506 1356 1509 1416
rect 1530 1373 1533 1526
rect 1554 1516 1557 1583
rect 1570 1536 1573 1616
rect 1570 1533 1589 1536
rect 1546 1513 1557 1516
rect 1546 1426 1549 1513
rect 1546 1423 1553 1426
rect 1538 1393 1541 1406
rect 1550 1356 1553 1423
rect 1562 1413 1565 1526
rect 1570 1513 1573 1526
rect 1594 1456 1597 1633
rect 1602 1603 1605 1616
rect 1610 1603 1613 1616
rect 1634 1613 1637 1633
rect 1666 1603 1669 1733
rect 1674 1603 1677 1806
rect 1714 1776 1717 1796
rect 1710 1773 1717 1776
rect 1682 1723 1685 1766
rect 1690 1696 1693 1726
rect 1682 1693 1693 1696
rect 1682 1596 1685 1693
rect 1674 1593 1685 1596
rect 1570 1453 1597 1456
rect 1562 1393 1565 1406
rect 1506 1353 1517 1356
rect 1498 1313 1501 1326
rect 1514 1306 1517 1353
rect 1510 1303 1517 1306
rect 1546 1353 1553 1356
rect 1466 1293 1477 1296
rect 1474 1236 1477 1293
rect 1466 1233 1477 1236
rect 1466 1213 1469 1233
rect 1458 1193 1461 1206
rect 1474 1123 1477 1166
rect 1458 1096 1461 1116
rect 1490 1113 1493 1206
rect 1498 1133 1501 1256
rect 1510 1246 1513 1303
rect 1546 1296 1549 1353
rect 1570 1316 1573 1453
rect 1586 1403 1589 1416
rect 1610 1393 1613 1416
rect 1618 1383 1621 1536
rect 1634 1456 1637 1586
rect 1650 1523 1653 1566
rect 1666 1516 1669 1526
rect 1642 1513 1669 1516
rect 1674 1513 1677 1593
rect 1698 1563 1701 1726
rect 1710 1706 1713 1773
rect 1722 1716 1725 1946
rect 1746 1803 1749 1926
rect 1802 1923 1805 1993
rect 1810 1933 1813 1986
rect 1818 1943 1821 2003
rect 1842 1983 1845 2016
rect 1858 2013 1861 2066
rect 1874 2016 1877 2113
rect 1906 2113 1917 2116
rect 1906 2046 1909 2113
rect 1906 2043 1917 2046
rect 1914 2026 1917 2043
rect 1866 2013 1877 2016
rect 1898 2023 1917 2026
rect 1898 2013 1901 2023
rect 1866 1956 1869 2013
rect 1866 1953 1873 1956
rect 1754 1736 1757 1816
rect 1738 1733 1757 1736
rect 1722 1713 1733 1716
rect 1710 1703 1717 1706
rect 1714 1553 1717 1703
rect 1714 1506 1717 1526
rect 1630 1453 1637 1456
rect 1706 1503 1717 1506
rect 1706 1456 1709 1503
rect 1706 1453 1717 1456
rect 1562 1313 1573 1316
rect 1594 1306 1597 1336
rect 1618 1316 1621 1376
rect 1630 1366 1633 1453
rect 1714 1433 1717 1453
rect 1630 1363 1637 1366
rect 1634 1343 1637 1363
rect 1666 1353 1669 1416
rect 1674 1403 1677 1426
rect 1706 1413 1709 1426
rect 1722 1416 1725 1526
rect 1730 1506 1733 1713
rect 1746 1713 1765 1716
rect 1738 1603 1741 1616
rect 1746 1613 1749 1713
rect 1754 1603 1757 1626
rect 1770 1613 1773 1916
rect 1850 1813 1853 1926
rect 1870 1906 1873 1953
rect 1882 1933 1885 1946
rect 1890 1926 1893 1996
rect 1906 1993 1909 2016
rect 1914 2013 1917 2023
rect 1922 2006 1925 2286
rect 1978 2236 1981 2446
rect 1986 2403 1989 2466
rect 1986 2333 1989 2376
rect 2002 2313 2005 2483
rect 2018 2403 2021 2526
rect 2050 2493 2053 2613
rect 2018 2393 2029 2396
rect 2034 2383 2037 2416
rect 2058 2403 2061 2606
rect 2070 2566 2073 2623
rect 2082 2576 2085 2873
rect 2106 2846 2109 2926
rect 2122 2913 2125 2936
rect 2138 2933 2141 2946
rect 2098 2843 2109 2846
rect 2090 2733 2093 2766
rect 2098 2733 2101 2843
rect 2106 2803 2109 2836
rect 2162 2826 2165 3040
rect 2170 2913 2173 2926
rect 2218 2923 2221 3040
rect 2322 2986 2325 3040
rect 2322 2983 2349 2986
rect 2290 2963 2333 2966
rect 2226 2943 2229 2956
rect 2290 2933 2293 2963
rect 2306 2933 2309 2946
rect 2282 2846 2285 2926
rect 2330 2923 2333 2963
rect 2346 2916 2349 2983
rect 2386 2923 2389 3040
rect 2402 2943 2405 2956
rect 2418 2926 2421 2946
rect 2410 2923 2421 2926
rect 2426 2923 2437 2926
rect 2338 2913 2349 2916
rect 2282 2843 2293 2846
rect 2162 2823 2173 2826
rect 2130 2803 2133 2816
rect 2154 2763 2157 2816
rect 2170 2746 2173 2823
rect 2210 2813 2213 2836
rect 2154 2743 2173 2746
rect 2090 2713 2101 2716
rect 2098 2686 2101 2713
rect 2098 2683 2117 2686
rect 2090 2596 2093 2626
rect 2098 2613 2101 2626
rect 2114 2613 2117 2683
rect 2122 2603 2125 2706
rect 2130 2603 2133 2636
rect 2090 2593 2141 2596
rect 2154 2586 2157 2743
rect 2162 2696 2165 2736
rect 2218 2733 2221 2816
rect 2234 2803 2237 2826
rect 2258 2803 2261 2816
rect 2290 2796 2293 2843
rect 2338 2836 2341 2913
rect 2410 2866 2413 2923
rect 2410 2863 2417 2866
rect 2330 2833 2341 2836
rect 2282 2793 2293 2796
rect 2178 2713 2181 2726
rect 2186 2713 2189 2726
rect 2162 2693 2181 2696
rect 2150 2583 2157 2586
rect 2082 2573 2117 2576
rect 2066 2563 2073 2566
rect 2066 2523 2069 2563
rect 2082 2533 2085 2546
rect 2114 2496 2117 2573
rect 2150 2526 2153 2583
rect 2178 2576 2181 2693
rect 2202 2613 2205 2716
rect 2242 2713 2245 2726
rect 2250 2706 2253 2726
rect 2218 2703 2253 2706
rect 2218 2616 2221 2703
rect 2226 2623 2245 2626
rect 2218 2613 2229 2616
rect 2242 2613 2245 2623
rect 2162 2573 2181 2576
rect 2098 2493 2117 2496
rect 2026 2323 2029 2376
rect 2074 2343 2077 2416
rect 2090 2343 2093 2366
rect 2098 2323 2101 2493
rect 2130 2486 2133 2526
rect 2150 2523 2157 2526
rect 2154 2506 2157 2523
rect 2162 2513 2165 2573
rect 2178 2533 2181 2546
rect 2154 2503 2165 2506
rect 2130 2483 2149 2486
rect 2138 2423 2141 2466
rect 2122 2413 2141 2416
rect 2114 2403 2133 2406
rect 2146 2403 2149 2483
rect 2162 2456 2165 2503
rect 2158 2453 2165 2456
rect 1930 2203 1933 2226
rect 1938 2203 1941 2236
rect 1946 2233 1981 2236
rect 1930 2123 1933 2196
rect 1914 2003 1925 2006
rect 1938 2106 1941 2136
rect 1946 2123 1949 2233
rect 1994 2203 1997 2226
rect 2002 2193 2005 2206
rect 1962 2143 1981 2146
rect 1954 2126 1957 2136
rect 1962 2133 1965 2143
rect 1954 2123 1965 2126
rect 1970 2106 1973 2136
rect 1938 2103 1973 2106
rect 1938 2003 1941 2103
rect 1978 2096 1981 2143
rect 1970 2093 1981 2096
rect 1898 1926 1901 1936
rect 1882 1923 1901 1926
rect 1914 1923 1917 2003
rect 1946 1986 1949 2046
rect 1938 1983 1949 1986
rect 1870 1903 1877 1906
rect 1874 1856 1877 1903
rect 1898 1883 1901 1916
rect 1866 1853 1877 1856
rect 1866 1833 1869 1853
rect 1786 1603 1789 1806
rect 1794 1763 1837 1766
rect 1794 1733 1797 1763
rect 1810 1733 1813 1746
rect 1834 1723 1837 1763
rect 1914 1756 1917 1816
rect 1922 1766 1925 1946
rect 1938 1856 1941 1983
rect 1938 1853 1945 1856
rect 1930 1823 1933 1836
rect 1942 1786 1945 1853
rect 1954 1833 1957 2016
rect 1970 2013 1973 2093
rect 1962 1993 1965 2006
rect 1978 1913 1981 1946
rect 1986 1856 1989 2016
rect 2002 1946 2005 2126
rect 2010 2123 2013 2216
rect 2018 2003 2021 2136
rect 2026 2123 2029 2276
rect 2106 2246 2109 2346
rect 2106 2243 2113 2246
rect 2034 2066 2037 2136
rect 2042 2123 2045 2196
rect 2050 2123 2053 2146
rect 2034 2063 2061 2066
rect 1994 1943 2005 1946
rect 1994 1933 1997 1943
rect 2026 1936 2029 1996
rect 2050 1936 2053 2016
rect 2058 2003 2061 2063
rect 2066 2013 2069 2216
rect 2082 2193 2085 2206
rect 2110 2176 2113 2243
rect 2122 2213 2125 2336
rect 2130 2323 2133 2403
rect 2158 2386 2161 2453
rect 2170 2426 2173 2446
rect 2210 2426 2213 2606
rect 2218 2573 2221 2606
rect 2274 2596 2277 2736
rect 2282 2733 2285 2793
rect 2306 2776 2309 2816
rect 2306 2773 2317 2776
rect 2314 2733 2317 2773
rect 2298 2713 2317 2716
rect 2298 2613 2301 2713
rect 2330 2656 2333 2833
rect 2338 2813 2341 2826
rect 2346 2733 2349 2816
rect 2362 2803 2365 2826
rect 2386 2803 2389 2816
rect 2402 2733 2405 2746
rect 2370 2713 2373 2726
rect 2378 2696 2381 2726
rect 2370 2693 2381 2696
rect 2330 2653 2341 2656
rect 2306 2603 2309 2616
rect 2314 2613 2317 2646
rect 2322 2613 2325 2626
rect 2338 2606 2341 2653
rect 2370 2626 2373 2693
rect 2414 2686 2417 2863
rect 2426 2743 2429 2923
rect 2442 2913 2445 2936
rect 2434 2736 2437 2816
rect 2466 2813 2469 2826
rect 2474 2796 2477 2946
rect 2498 2913 2501 2926
rect 2554 2923 2557 3040
rect 2578 2933 2581 2946
rect 2466 2793 2477 2796
rect 2434 2733 2445 2736
rect 2426 2706 2429 2726
rect 2426 2703 2433 2706
rect 2414 2683 2421 2686
rect 2370 2623 2381 2626
rect 2330 2603 2341 2606
rect 2378 2606 2381 2623
rect 2386 2613 2389 2676
rect 2402 2613 2405 2656
rect 2378 2603 2389 2606
rect 2266 2593 2277 2596
rect 2266 2533 2269 2593
rect 2306 2533 2309 2546
rect 2226 2436 2229 2526
rect 2226 2433 2237 2436
rect 2170 2423 2181 2426
rect 2154 2383 2161 2386
rect 2138 2256 2141 2326
rect 2154 2276 2157 2383
rect 2178 2376 2181 2423
rect 2170 2373 2181 2376
rect 2170 2286 2173 2373
rect 2170 2283 2181 2286
rect 2154 2273 2165 2276
rect 2138 2253 2153 2256
rect 2150 2206 2153 2253
rect 2162 2213 2165 2273
rect 2178 2206 2181 2283
rect 2150 2203 2157 2206
rect 2106 2173 2113 2176
rect 2106 2156 2109 2173
rect 2090 2153 2109 2156
rect 2090 1966 2093 2153
rect 2114 2133 2117 2146
rect 2130 2133 2133 2196
rect 2114 2013 2117 2126
rect 2090 1963 2109 1966
rect 2026 1933 2033 1936
rect 2018 1883 2021 1926
rect 1986 1853 2021 1856
rect 1942 1783 1949 1786
rect 1922 1763 1941 1766
rect 1898 1753 1917 1756
rect 1890 1703 1893 1726
rect 1898 1713 1901 1753
rect 1914 1733 1917 1746
rect 1938 1676 1941 1763
rect 1946 1703 1949 1783
rect 1930 1673 1941 1676
rect 1738 1533 1741 1546
rect 1754 1506 1757 1536
rect 1730 1503 1757 1506
rect 1722 1413 1733 1416
rect 1674 1333 1677 1396
rect 1722 1383 1725 1406
rect 1570 1303 1597 1306
rect 1610 1313 1621 1316
rect 1546 1293 1557 1296
rect 1506 1243 1513 1246
rect 1506 1176 1509 1243
rect 1506 1173 1513 1176
rect 1510 1106 1513 1173
rect 1458 1093 1469 1096
rect 1466 1036 1469 1093
rect 1482 1056 1485 1106
rect 1506 1103 1513 1106
rect 1506 1083 1509 1103
rect 1482 1053 1493 1056
rect 1462 1033 1469 1036
rect 1490 1036 1493 1053
rect 1490 1033 1497 1036
rect 1462 976 1465 1033
rect 1474 993 1477 1016
rect 1494 976 1497 1033
rect 1506 1003 1509 1016
rect 1434 943 1453 946
rect 1458 973 1465 976
rect 1490 973 1497 976
rect 1434 653 1437 943
rect 1442 813 1445 936
rect 1458 883 1461 973
rect 1466 933 1469 956
rect 1490 926 1493 973
rect 1514 963 1517 1016
rect 1522 986 1525 1206
rect 1554 1186 1557 1293
rect 1610 1236 1613 1313
rect 1674 1306 1677 1326
rect 1698 1306 1701 1326
rect 1610 1233 1621 1236
rect 1546 1183 1557 1186
rect 1546 1116 1549 1183
rect 1562 1143 1565 1216
rect 1602 1166 1605 1216
rect 1594 1163 1605 1166
rect 1610 1163 1613 1206
rect 1530 1096 1533 1116
rect 1546 1113 1557 1116
rect 1562 1113 1565 1126
rect 1530 1093 1541 1096
rect 1538 1026 1541 1093
rect 1530 1023 1541 1026
rect 1530 1003 1533 1023
rect 1554 1016 1557 1113
rect 1594 1086 1597 1163
rect 1610 1096 1613 1136
rect 1618 1123 1621 1233
rect 1626 1193 1629 1306
rect 1674 1303 1701 1306
rect 1682 1243 1717 1246
rect 1650 1223 1653 1236
rect 1682 1223 1685 1243
rect 1698 1223 1701 1236
rect 1714 1223 1717 1243
rect 1722 1216 1725 1326
rect 1698 1213 1725 1216
rect 1730 1196 1733 1413
rect 1738 1386 1741 1436
rect 1746 1403 1749 1503
rect 1794 1486 1797 1526
rect 1786 1483 1797 1486
rect 1786 1426 1789 1483
rect 1754 1393 1757 1406
rect 1738 1383 1745 1386
rect 1742 1226 1745 1383
rect 1610 1093 1621 1096
rect 1594 1083 1605 1086
rect 1602 1063 1605 1083
rect 1618 1026 1621 1093
rect 1610 1023 1621 1026
rect 1554 1013 1565 1016
rect 1554 993 1557 1006
rect 1522 983 1549 986
rect 1474 903 1477 926
rect 1486 923 1493 926
rect 1486 876 1489 923
rect 1498 883 1501 916
rect 1514 896 1517 946
rect 1522 926 1525 976
rect 1546 933 1549 983
rect 1522 923 1557 926
rect 1562 923 1565 1013
rect 1586 983 1589 1006
rect 1610 976 1613 1023
rect 1634 1013 1637 1136
rect 1650 1106 1653 1126
rect 1690 1123 1693 1196
rect 1722 1193 1733 1196
rect 1738 1223 1745 1226
rect 1706 1116 1709 1126
rect 1682 1113 1709 1116
rect 1650 1103 1661 1106
rect 1658 1016 1661 1103
rect 1722 1096 1725 1193
rect 1738 1103 1741 1223
rect 1746 1183 1749 1206
rect 1754 1133 1757 1376
rect 1762 1333 1765 1426
rect 1786 1423 1797 1426
rect 1794 1403 1797 1423
rect 1770 1333 1773 1356
rect 1786 1333 1789 1376
rect 1762 1323 1773 1326
rect 1770 1286 1773 1323
rect 1778 1303 1781 1326
rect 1770 1283 1781 1286
rect 1778 1236 1781 1283
rect 1770 1233 1781 1236
rect 1770 1193 1773 1233
rect 1802 1163 1805 1616
rect 1850 1603 1853 1616
rect 1858 1593 1861 1616
rect 1858 1556 1861 1586
rect 1842 1553 1861 1556
rect 1810 1393 1813 1406
rect 1826 1333 1829 1416
rect 1842 1403 1845 1553
rect 1850 1513 1853 1526
rect 1866 1463 1869 1536
rect 1890 1523 1893 1606
rect 1898 1603 1901 1616
rect 1930 1576 1933 1673
rect 1930 1573 1937 1576
rect 1934 1496 1937 1573
rect 1946 1506 1949 1696
rect 1954 1683 1957 1826
rect 1994 1773 1997 1806
rect 2018 1796 2021 1853
rect 2010 1793 2021 1796
rect 2010 1756 2013 1793
rect 2030 1776 2033 1933
rect 2042 1813 2045 1936
rect 2050 1933 2069 1936
rect 2090 1933 2093 1946
rect 2066 1916 2069 1933
rect 2066 1913 2077 1916
rect 2006 1753 2013 1756
rect 2026 1773 2033 1776
rect 1962 1613 1965 1726
rect 1978 1606 1981 1746
rect 1994 1623 1997 1726
rect 2006 1636 2009 1753
rect 2026 1733 2029 1773
rect 2058 1766 2061 1886
rect 2074 1776 2077 1913
rect 2098 1853 2101 1926
rect 2106 1896 2109 1963
rect 2122 1933 2125 1996
rect 2138 1946 2141 2076
rect 2154 1956 2157 2203
rect 2170 2203 2181 2206
rect 2170 2156 2173 2203
rect 2170 2153 2177 2156
rect 2162 2123 2165 2146
rect 2174 2106 2177 2153
rect 2170 2103 2177 2106
rect 2170 2083 2173 2103
rect 2194 2073 2197 2416
rect 2202 2403 2205 2426
rect 2210 2423 2221 2426
rect 2218 2406 2221 2423
rect 2210 2403 2221 2406
rect 2234 2403 2237 2433
rect 2258 2423 2261 2446
rect 2282 2413 2285 2526
rect 2330 2496 2333 2603
rect 2322 2493 2333 2496
rect 2322 2436 2325 2493
rect 2314 2433 2325 2436
rect 2202 2213 2205 2226
rect 2210 2213 2213 2403
rect 2266 2383 2269 2396
rect 2226 2333 2229 2356
rect 2218 2223 2221 2236
rect 2202 2123 2213 2126
rect 2218 2113 2221 2126
rect 2162 2023 2165 2046
rect 2186 2003 2189 2026
rect 2202 1993 2205 2006
rect 2154 1953 2161 1956
rect 2138 1943 2149 1946
rect 2106 1893 2113 1896
rect 2054 1763 2061 1766
rect 2066 1773 2077 1776
rect 2006 1633 2013 1636
rect 1970 1603 1981 1606
rect 1970 1533 1973 1603
rect 1986 1583 1989 1616
rect 2002 1603 2005 1616
rect 2010 1586 2013 1633
rect 2018 1593 2021 1706
rect 2054 1686 2057 1763
rect 2066 1696 2069 1773
rect 2090 1753 2093 1816
rect 2074 1723 2077 1736
rect 2066 1693 2073 1696
rect 2042 1666 2045 1686
rect 2054 1683 2061 1686
rect 2034 1663 2045 1666
rect 2034 1596 2037 1663
rect 2050 1603 2053 1666
rect 2034 1593 2045 1596
rect 2002 1583 2013 1586
rect 1954 1513 1957 1526
rect 2002 1516 2005 1583
rect 2018 1523 2021 1556
rect 2042 1536 2045 1593
rect 2038 1533 2045 1536
rect 2002 1513 2013 1516
rect 1946 1503 1965 1506
rect 1934 1493 1941 1496
rect 1762 1106 1765 1136
rect 1810 1133 1813 1196
rect 1818 1123 1821 1236
rect 1834 1226 1837 1326
rect 1858 1303 1861 1316
rect 1874 1306 1877 1406
rect 1898 1366 1901 1416
rect 1938 1413 1941 1493
rect 1954 1393 1957 1416
rect 1882 1363 1901 1366
rect 1882 1333 1885 1363
rect 1898 1306 1901 1336
rect 1946 1323 1949 1336
rect 1874 1303 1901 1306
rect 1962 1276 1965 1503
rect 1954 1273 1965 1276
rect 1834 1223 1853 1226
rect 1762 1103 1797 1106
rect 1722 1093 1733 1096
rect 1650 1013 1661 1016
rect 1594 973 1613 976
rect 1514 893 1533 896
rect 1486 873 1493 876
rect 1450 736 1453 836
rect 1490 826 1493 873
rect 1490 823 1501 826
rect 1474 813 1493 816
rect 1498 776 1501 823
rect 1514 793 1517 806
rect 1498 773 1509 776
rect 1442 733 1453 736
rect 1458 763 1501 766
rect 1458 733 1461 763
rect 1474 733 1477 746
rect 1442 696 1445 733
rect 1450 713 1453 726
rect 1498 723 1501 763
rect 1442 693 1453 696
rect 1506 693 1509 773
rect 1530 766 1533 893
rect 1578 836 1581 936
rect 1594 933 1597 973
rect 1650 933 1653 1013
rect 1626 853 1629 926
rect 1570 833 1581 836
rect 1554 793 1557 816
rect 1522 763 1533 766
rect 1434 613 1437 626
rect 1450 616 1453 693
rect 1450 613 1469 616
rect 1482 613 1485 636
rect 1442 593 1445 606
rect 1434 533 1437 546
rect 1466 543 1469 613
rect 1506 603 1509 626
rect 1522 566 1525 763
rect 1570 733 1573 833
rect 1618 796 1621 816
rect 1634 803 1637 906
rect 1610 793 1621 796
rect 1610 746 1613 793
rect 1610 743 1621 746
rect 1666 743 1669 956
rect 1682 813 1685 936
rect 1698 923 1701 1016
rect 1706 893 1709 1016
rect 1714 986 1717 1066
rect 1730 1016 1733 1093
rect 1722 1013 1733 1016
rect 1722 1003 1725 1013
rect 1714 983 1721 986
rect 1718 886 1721 983
rect 1746 976 1749 1006
rect 1770 996 1773 1016
rect 1714 883 1721 886
rect 1738 973 1749 976
rect 1714 826 1717 883
rect 1738 843 1741 973
rect 1754 953 1757 996
rect 1766 993 1773 996
rect 1766 866 1769 993
rect 1778 923 1781 1006
rect 1786 916 1789 1036
rect 1794 1013 1797 1103
rect 1818 1003 1821 1026
rect 1826 1013 1829 1136
rect 1834 1123 1837 1223
rect 1842 1116 1845 1216
rect 1850 1203 1853 1223
rect 1858 1216 1861 1236
rect 1858 1213 1869 1216
rect 1858 1173 1861 1206
rect 1850 1123 1853 1166
rect 1842 1113 1853 1116
rect 1866 1073 1869 1213
rect 1954 1186 1957 1273
rect 1970 1263 1973 1416
rect 1978 1326 1981 1356
rect 2010 1346 2013 1513
rect 2038 1426 2041 1533
rect 2018 1413 2021 1426
rect 2038 1423 2045 1426
rect 2034 1346 2037 1406
rect 1994 1343 2037 1346
rect 1978 1323 1989 1326
rect 1994 1216 1997 1343
rect 2002 1316 2005 1336
rect 2018 1333 2029 1336
rect 2018 1323 2029 1326
rect 2034 1323 2037 1336
rect 2018 1316 2021 1323
rect 2042 1316 2045 1423
rect 2050 1373 2053 1526
rect 2058 1493 2061 1683
rect 2070 1506 2073 1693
rect 2098 1676 2101 1846
rect 2110 1826 2113 1893
rect 2106 1823 2113 1826
rect 2106 1786 2109 1823
rect 2114 1793 2117 1806
rect 2122 1803 2125 1856
rect 2146 1786 2149 1943
rect 2158 1906 2161 1953
rect 2154 1903 2161 1906
rect 2154 1843 2157 1903
rect 2162 1823 2165 1886
rect 2170 1803 2173 1926
rect 2202 1923 2205 1946
rect 2226 1906 2229 2226
rect 2234 2203 2237 2216
rect 2242 2196 2245 2346
rect 2274 2323 2277 2406
rect 2290 2403 2293 2416
rect 2314 2376 2317 2433
rect 2330 2403 2333 2426
rect 2346 2416 2349 2526
rect 2386 2523 2389 2603
rect 2394 2593 2397 2606
rect 2402 2506 2405 2606
rect 2410 2593 2413 2666
rect 2394 2503 2405 2506
rect 2346 2413 2357 2416
rect 2354 2403 2357 2413
rect 2314 2373 2325 2376
rect 2322 2323 2325 2373
rect 2362 2366 2365 2426
rect 2394 2416 2397 2503
rect 2394 2413 2405 2416
rect 2410 2413 2413 2526
rect 2418 2496 2421 2683
rect 2430 2636 2433 2703
rect 2442 2673 2445 2716
rect 2426 2633 2433 2636
rect 2426 2613 2429 2633
rect 2466 2576 2469 2793
rect 2466 2573 2477 2576
rect 2418 2493 2429 2496
rect 2338 2363 2365 2366
rect 2338 2273 2341 2363
rect 2354 2333 2357 2346
rect 2378 2323 2381 2396
rect 2394 2383 2397 2396
rect 2234 2193 2245 2196
rect 2282 2136 2285 2146
rect 2234 2133 2285 2136
rect 2290 2133 2293 2196
rect 2234 2013 2237 2026
rect 2218 1903 2229 1906
rect 2106 1783 2133 1786
rect 2114 1716 2117 1736
rect 2090 1673 2101 1676
rect 2110 1713 2117 1716
rect 2090 1626 2093 1673
rect 2110 1636 2113 1713
rect 2122 1663 2125 1726
rect 2082 1623 2093 1626
rect 2106 1633 2113 1636
rect 2082 1546 2085 1623
rect 2106 1616 2109 1633
rect 2090 1613 2109 1616
rect 2090 1593 2093 1606
rect 2082 1543 2101 1546
rect 2066 1503 2073 1506
rect 2066 1486 2069 1503
rect 2062 1483 2069 1486
rect 2062 1386 2065 1483
rect 2074 1396 2077 1466
rect 2082 1413 2085 1536
rect 2090 1503 2093 1526
rect 2098 1486 2101 1543
rect 2106 1533 2109 1556
rect 2106 1493 2109 1516
rect 2094 1483 2101 1486
rect 2074 1393 2085 1396
rect 2062 1383 2069 1386
rect 2002 1313 2021 1316
rect 2026 1313 2061 1316
rect 2050 1223 2053 1306
rect 1978 1213 1997 1216
rect 1954 1183 1961 1186
rect 1874 1096 1877 1136
rect 1874 1093 1881 1096
rect 1878 1036 1881 1093
rect 1874 1033 1881 1036
rect 1874 1013 1877 1033
rect 1850 986 1853 1006
rect 1802 983 1853 986
rect 1778 913 1789 916
rect 1766 863 1773 866
rect 1706 823 1717 826
rect 1546 613 1549 626
rect 1522 563 1533 566
rect 1426 523 1445 526
rect 1426 483 1429 516
rect 1442 456 1445 523
rect 1490 503 1493 526
rect 1434 453 1445 456
rect 1330 383 1381 386
rect 1282 313 1293 316
rect 1298 296 1301 336
rect 1290 293 1301 296
rect 1290 236 1293 293
rect 1314 243 1317 336
rect 1370 333 1373 356
rect 1378 256 1381 383
rect 1370 253 1381 256
rect 1402 253 1405 403
rect 1426 373 1429 416
rect 1410 323 1413 336
rect 1434 326 1437 453
rect 1442 413 1445 436
rect 1442 383 1445 406
rect 1418 323 1437 326
rect 1442 313 1445 376
rect 1450 256 1453 336
rect 1474 323 1477 416
rect 1490 413 1493 426
rect 1498 406 1501 546
rect 1506 466 1509 536
rect 1514 486 1517 536
rect 1530 533 1533 563
rect 1554 533 1557 726
rect 1610 713 1613 726
rect 1602 566 1605 616
rect 1610 583 1613 596
rect 1570 563 1605 566
rect 1570 546 1573 563
rect 1566 543 1573 546
rect 1554 486 1557 526
rect 1514 483 1557 486
rect 1506 463 1513 466
rect 1490 403 1501 406
rect 1490 356 1493 403
rect 1510 396 1513 463
rect 1566 436 1569 543
rect 1566 433 1573 436
rect 1486 353 1493 356
rect 1506 393 1513 396
rect 1522 413 1549 416
rect 1486 306 1489 353
rect 1434 253 1453 256
rect 1482 303 1489 306
rect 1290 233 1301 236
rect 1298 213 1301 233
rect 1330 213 1333 226
rect 1370 216 1373 253
rect 1354 213 1373 216
rect 1434 213 1437 253
rect 1482 236 1485 303
rect 1482 233 1493 236
rect 1250 193 1253 206
rect 1298 163 1341 166
rect 1250 133 1253 146
rect 1298 123 1301 163
rect 1338 133 1341 163
rect 1346 143 1349 156
rect 1354 126 1357 213
rect 1362 203 1373 206
rect 1386 193 1389 206
rect 1474 203 1477 216
rect 1490 176 1493 233
rect 1458 173 1493 176
rect 1498 173 1501 346
rect 1506 323 1509 393
rect 1522 313 1525 413
rect 1538 356 1541 406
rect 1554 393 1557 406
rect 1562 403 1565 416
rect 1570 373 1573 433
rect 1578 356 1581 556
rect 1618 546 1621 743
rect 1650 626 1653 726
rect 1658 723 1661 736
rect 1610 543 1621 546
rect 1630 623 1653 626
rect 1610 466 1613 543
rect 1630 536 1633 623
rect 1642 613 1653 616
rect 1642 546 1645 613
rect 1650 576 1653 606
rect 1666 593 1669 606
rect 1690 576 1693 616
rect 1650 573 1693 576
rect 1642 543 1653 546
rect 1630 533 1637 536
rect 1610 463 1621 466
rect 1538 353 1589 356
rect 1538 333 1541 346
rect 1586 333 1589 353
rect 1594 343 1597 406
rect 1618 386 1621 463
rect 1614 383 1621 386
rect 1538 276 1541 326
rect 1538 273 1557 276
rect 1554 213 1557 273
rect 1562 206 1565 326
rect 1570 306 1573 326
rect 1594 323 1597 336
rect 1594 306 1597 316
rect 1570 303 1597 306
rect 1506 203 1517 206
rect 1530 193 1533 206
rect 1558 203 1565 206
rect 1426 133 1429 146
rect 1138 63 1149 66
rect 1138 0 1141 63
rect 1154 0 1157 56
rect 1330 0 1333 126
rect 1354 123 1381 126
rect 1458 116 1461 173
rect 1474 163 1493 166
rect 1474 123 1477 163
rect 1490 136 1493 163
rect 1506 143 1517 146
rect 1490 133 1517 136
rect 1458 113 1469 116
rect 1466 93 1469 113
rect 1506 0 1509 126
rect 1546 123 1549 176
rect 1558 126 1561 203
rect 1554 123 1561 126
rect 1554 106 1557 123
rect 1546 103 1557 106
rect 1546 16 1549 103
rect 1546 13 1557 16
rect 1554 0 1557 13
rect 1570 0 1573 256
rect 1602 196 1605 376
rect 1614 326 1617 383
rect 1614 323 1621 326
rect 1610 293 1613 306
rect 1610 203 1613 216
rect 1602 193 1613 196
rect 1586 133 1589 146
rect 1586 0 1589 126
rect 1610 123 1613 193
rect 1602 0 1605 96
rect 1618 0 1621 323
rect 1626 76 1629 526
rect 1634 396 1637 533
rect 1642 506 1645 536
rect 1650 523 1653 543
rect 1682 523 1685 566
rect 1698 553 1701 736
rect 1706 543 1709 823
rect 1714 566 1717 816
rect 1762 813 1765 846
rect 1770 806 1773 863
rect 1778 823 1781 913
rect 1722 723 1725 806
rect 1762 803 1773 806
rect 1738 733 1741 786
rect 1762 746 1765 803
rect 1762 743 1769 746
rect 1766 696 1769 743
rect 1778 723 1781 806
rect 1762 693 1769 696
rect 1714 563 1725 566
rect 1698 526 1701 536
rect 1690 523 1701 526
rect 1642 503 1677 506
rect 1642 413 1645 466
rect 1634 393 1641 396
rect 1638 246 1641 393
rect 1634 243 1641 246
rect 1634 186 1637 243
rect 1650 193 1653 346
rect 1658 323 1661 396
rect 1666 313 1669 376
rect 1674 353 1677 503
rect 1690 463 1693 523
rect 1722 516 1725 563
rect 1714 513 1725 516
rect 1714 426 1717 513
rect 1690 413 1693 426
rect 1698 423 1717 426
rect 1674 323 1677 336
rect 1634 183 1653 186
rect 1650 166 1653 183
rect 1650 163 1657 166
rect 1634 123 1637 136
rect 1654 86 1657 163
rect 1674 143 1677 156
rect 1666 133 1677 136
rect 1666 106 1669 126
rect 1682 123 1685 396
rect 1690 333 1693 406
rect 1698 346 1701 423
rect 1706 353 1709 416
rect 1714 413 1725 416
rect 1714 363 1717 406
rect 1730 373 1733 396
rect 1746 393 1749 616
rect 1762 533 1765 693
rect 1802 686 1805 776
rect 1810 696 1813 983
rect 1850 976 1853 983
rect 1890 976 1893 1136
rect 1938 1123 1941 1166
rect 1958 1116 1961 1183
rect 1970 1123 1973 1176
rect 1958 1113 1965 1116
rect 1962 1093 1965 1113
rect 1978 1036 1981 1213
rect 1986 1203 1997 1206
rect 1994 1186 1997 1203
rect 1994 1183 2013 1186
rect 1986 1096 1989 1176
rect 2010 1123 2013 1183
rect 2018 1163 2021 1206
rect 2018 1133 2021 1146
rect 2034 1106 2037 1166
rect 2018 1103 2037 1106
rect 1986 1093 1997 1096
rect 1970 1033 1981 1036
rect 1930 1013 1933 1026
rect 1946 993 1949 1006
rect 1850 973 1893 976
rect 1858 943 1901 946
rect 1858 933 1861 943
rect 1882 926 1885 936
rect 1834 826 1837 926
rect 1842 843 1845 926
rect 1874 923 1885 926
rect 1874 916 1877 923
rect 1866 913 1877 916
rect 1890 913 1893 926
rect 1866 866 1869 913
rect 1858 863 1869 866
rect 1834 823 1841 826
rect 1838 766 1841 823
rect 1858 813 1861 863
rect 1890 806 1893 816
rect 1898 813 1901 943
rect 1930 933 1933 986
rect 1962 913 1965 926
rect 1970 923 1973 1033
rect 1986 933 1989 1016
rect 1954 853 1973 856
rect 1954 813 1957 853
rect 1890 803 1901 806
rect 1898 766 1901 803
rect 1962 796 1965 846
rect 1970 813 1973 853
rect 1838 763 1877 766
rect 1898 763 1909 766
rect 1834 733 1837 746
rect 1818 713 1821 726
rect 1866 706 1869 726
rect 1862 703 1869 706
rect 1810 693 1821 696
rect 1802 683 1813 686
rect 1770 603 1773 616
rect 1802 613 1805 626
rect 1770 533 1773 546
rect 1778 523 1781 606
rect 1810 593 1813 683
rect 1818 586 1821 693
rect 1810 583 1821 586
rect 1810 533 1813 583
rect 1754 513 1765 516
rect 1778 413 1789 416
rect 1698 343 1717 346
rect 1698 333 1709 336
rect 1698 213 1701 333
rect 1714 256 1717 343
rect 1722 313 1725 356
rect 1778 353 1781 413
rect 1794 403 1797 426
rect 1802 396 1805 416
rect 1834 413 1837 696
rect 1862 636 1865 703
rect 1862 633 1869 636
rect 1842 603 1853 606
rect 1786 393 1805 396
rect 1714 253 1721 256
rect 1718 186 1721 253
rect 1714 183 1721 186
rect 1730 216 1733 336
rect 1778 323 1781 336
rect 1786 333 1789 376
rect 1842 336 1845 546
rect 1850 523 1853 603
rect 1858 593 1861 616
rect 1866 603 1869 633
rect 1874 456 1877 763
rect 1882 516 1885 756
rect 1906 686 1909 763
rect 1954 753 1957 796
rect 1962 793 1973 796
rect 1898 683 1909 686
rect 1898 643 1901 683
rect 1898 553 1901 616
rect 1922 556 1925 736
rect 1962 733 1965 746
rect 1930 706 1933 726
rect 1970 723 1973 793
rect 1994 743 1997 1093
rect 2018 1026 2021 1103
rect 2014 1023 2021 1026
rect 2014 966 2017 1023
rect 2026 983 2029 1016
rect 2034 973 2037 1016
rect 2014 963 2021 966
rect 2002 776 2005 806
rect 2018 803 2021 963
rect 2026 903 2029 916
rect 2050 913 2053 926
rect 2058 823 2061 1313
rect 2066 1303 2069 1383
rect 2082 1296 2085 1393
rect 2074 1293 2085 1296
rect 2074 1163 2077 1293
rect 2094 1256 2097 1483
rect 2094 1253 2101 1256
rect 2098 1176 2101 1253
rect 2082 1173 2101 1176
rect 2106 1173 2109 1476
rect 2114 1426 2117 1526
rect 2130 1503 2133 1783
rect 2138 1783 2149 1786
rect 2138 1643 2141 1783
rect 2146 1726 2149 1776
rect 2154 1733 2165 1736
rect 2146 1723 2157 1726
rect 2138 1576 2141 1606
rect 2154 1603 2157 1723
rect 2186 1673 2189 1836
rect 2218 1816 2221 1903
rect 2234 1826 2237 1926
rect 2250 1893 2253 1926
rect 2234 1823 2253 1826
rect 2210 1813 2221 1816
rect 2234 1813 2245 1816
rect 2250 1813 2253 1823
rect 2258 1813 2261 1956
rect 2266 1906 2269 2116
rect 2274 1923 2277 2076
rect 2282 2026 2285 2133
rect 2290 2063 2293 2126
rect 2306 2113 2309 2216
rect 2354 2203 2357 2246
rect 2402 2243 2405 2413
rect 2426 2406 2429 2493
rect 2418 2403 2429 2406
rect 2418 2366 2421 2403
rect 2418 2363 2429 2366
rect 2426 2286 2429 2363
rect 2410 2283 2429 2286
rect 2410 2236 2413 2283
rect 2442 2256 2445 2546
rect 2474 2536 2477 2573
rect 2490 2543 2493 2816
rect 2506 2733 2517 2736
rect 2530 2733 2533 2816
rect 2570 2813 2597 2816
rect 2570 2733 2573 2813
rect 2610 2803 2613 2926
rect 2658 2923 2661 3040
rect 2762 2976 2765 3040
rect 2762 2973 2773 2976
rect 2682 2933 2685 2946
rect 2618 2813 2637 2816
rect 2698 2813 2709 2816
rect 2618 2793 2637 2796
rect 2634 2773 2637 2793
rect 2698 2776 2701 2813
rect 2714 2803 2717 2926
rect 2770 2923 2773 2973
rect 2786 2933 2789 2946
rect 2834 2866 2837 2926
rect 2866 2923 2869 3040
rect 2834 2863 2861 2866
rect 2722 2793 2725 2806
rect 2690 2773 2701 2776
rect 2514 2726 2517 2733
rect 2506 2653 2509 2726
rect 2514 2723 2533 2726
rect 2522 2713 2533 2716
rect 2498 2613 2501 2626
rect 2506 2603 2509 2616
rect 2522 2613 2525 2713
rect 2514 2603 2525 2606
rect 2466 2533 2477 2536
rect 2466 2416 2469 2533
rect 2458 2413 2469 2416
rect 2474 2413 2477 2426
rect 2482 2416 2485 2526
rect 2522 2523 2525 2603
rect 2530 2506 2533 2656
rect 2538 2616 2541 2636
rect 2538 2613 2557 2616
rect 2578 2613 2581 2656
rect 2538 2573 2541 2606
rect 2522 2503 2533 2506
rect 2498 2423 2501 2466
rect 2522 2416 2525 2503
rect 2482 2413 2493 2416
rect 2522 2413 2533 2416
rect 2458 2353 2461 2413
rect 2466 2403 2477 2406
rect 2490 2403 2493 2413
rect 2458 2293 2461 2326
rect 2474 2303 2477 2396
rect 2498 2323 2501 2396
rect 2514 2363 2517 2396
rect 2530 2366 2533 2413
rect 2538 2403 2541 2526
rect 2554 2496 2557 2613
rect 2594 2603 2597 2616
rect 2618 2583 2621 2736
rect 2634 2733 2637 2746
rect 2634 2633 2637 2726
rect 2626 2613 2629 2626
rect 2642 2623 2653 2626
rect 2658 2616 2661 2726
rect 2682 2696 2685 2736
rect 2690 2733 2693 2773
rect 2674 2693 2685 2696
rect 2634 2613 2661 2616
rect 2658 2596 2661 2606
rect 2666 2603 2669 2616
rect 2674 2596 2677 2693
rect 2690 2606 2693 2726
rect 2714 2613 2717 2706
rect 2754 2703 2757 2716
rect 2690 2603 2725 2606
rect 2658 2593 2677 2596
rect 2578 2533 2581 2546
rect 2658 2526 2661 2593
rect 2730 2566 2733 2646
rect 2738 2603 2741 2616
rect 2730 2563 2749 2566
rect 2674 2533 2677 2546
rect 2554 2493 2565 2496
rect 2546 2413 2549 2426
rect 2562 2376 2565 2493
rect 2610 2416 2613 2426
rect 2618 2423 2621 2446
rect 2610 2413 2621 2416
rect 2610 2406 2613 2413
rect 2594 2403 2613 2406
rect 2626 2403 2629 2526
rect 2650 2523 2661 2526
rect 2650 2403 2653 2523
rect 2722 2506 2725 2526
rect 2714 2503 2725 2506
rect 2666 2413 2669 2436
rect 2690 2403 2693 2496
rect 2714 2446 2717 2503
rect 2746 2486 2749 2563
rect 2738 2483 2749 2486
rect 2714 2443 2725 2446
rect 2522 2363 2533 2366
rect 2546 2373 2565 2376
rect 2714 2373 2717 2426
rect 2722 2403 2725 2443
rect 2722 2383 2725 2396
rect 2738 2376 2741 2483
rect 2762 2466 2765 2806
rect 2770 2653 2773 2726
rect 2778 2716 2781 2776
rect 2794 2733 2797 2816
rect 2842 2793 2845 2816
rect 2858 2803 2861 2863
rect 2850 2773 2853 2796
rect 2890 2766 2893 2816
rect 2874 2763 2893 2766
rect 2802 2733 2829 2736
rect 2850 2733 2853 2746
rect 2826 2726 2829 2733
rect 2826 2723 2837 2726
rect 2778 2713 2789 2716
rect 2786 2646 2789 2713
rect 2778 2643 2789 2646
rect 2802 2713 2829 2716
rect 2778 2486 2781 2643
rect 2802 2613 2805 2713
rect 2794 2533 2797 2606
rect 2802 2493 2805 2526
rect 2810 2486 2813 2546
rect 2754 2463 2765 2466
rect 2770 2483 2813 2486
rect 2754 2396 2757 2463
rect 2754 2393 2765 2396
rect 2770 2393 2773 2483
rect 2778 2416 2781 2426
rect 2778 2413 2789 2416
rect 2794 2403 2797 2426
rect 2762 2376 2765 2393
rect 2738 2373 2749 2376
rect 2762 2373 2781 2376
rect 2522 2323 2525 2363
rect 2546 2356 2549 2373
rect 2542 2353 2549 2356
rect 2402 2233 2413 2236
rect 2418 2253 2445 2256
rect 2542 2256 2545 2353
rect 2554 2266 2557 2366
rect 2626 2363 2645 2366
rect 2578 2333 2581 2356
rect 2562 2313 2565 2326
rect 2626 2323 2629 2363
rect 2642 2336 2645 2363
rect 2642 2333 2669 2336
rect 2674 2323 2677 2346
rect 2682 2276 2685 2346
rect 2730 2333 2733 2366
rect 2746 2326 2749 2373
rect 2666 2273 2685 2276
rect 2554 2263 2561 2266
rect 2542 2253 2549 2256
rect 2362 2153 2365 2216
rect 2378 2213 2381 2226
rect 2402 2186 2405 2233
rect 2418 2203 2421 2253
rect 2402 2183 2413 2186
rect 2330 2113 2333 2136
rect 2378 2133 2381 2146
rect 2354 2106 2357 2126
rect 2298 2103 2357 2106
rect 2282 2023 2301 2026
rect 2282 2013 2285 2023
rect 2266 1903 2277 1906
rect 2210 1666 2213 1813
rect 2274 1806 2277 1903
rect 2290 1813 2293 2016
rect 2298 2003 2301 2023
rect 2338 2013 2341 2036
rect 2306 1933 2309 1966
rect 2354 1943 2357 2086
rect 2226 1793 2229 1806
rect 2234 1803 2277 1806
rect 2226 1746 2229 1766
rect 2222 1743 2229 1746
rect 2222 1696 2225 1743
rect 2234 1703 2237 1803
rect 2242 1696 2245 1736
rect 2266 1703 2269 1726
rect 2274 1696 2277 1726
rect 2222 1693 2229 1696
rect 2242 1693 2277 1696
rect 2226 1676 2229 1693
rect 2226 1673 2233 1676
rect 2210 1663 2221 1666
rect 2202 1613 2205 1626
rect 2138 1573 2205 1576
rect 2218 1573 2221 1663
rect 2230 1576 2233 1673
rect 2242 1603 2245 1626
rect 2266 1613 2269 1626
rect 2226 1573 2233 1576
rect 2250 1576 2253 1606
rect 2290 1603 2293 1806
rect 2306 1746 2309 1926
rect 2354 1923 2357 1936
rect 2362 1923 2365 2066
rect 2410 2056 2413 2183
rect 2426 2103 2429 2136
rect 2442 2133 2445 2206
rect 2458 2166 2461 2216
rect 2498 2203 2501 2216
rect 2522 2166 2525 2206
rect 2546 2196 2549 2253
rect 2454 2163 2461 2166
rect 2490 2163 2525 2166
rect 2538 2193 2549 2196
rect 2402 2053 2413 2056
rect 2370 1933 2373 1966
rect 2346 1846 2349 1856
rect 2322 1843 2349 1846
rect 2322 1763 2325 1843
rect 2330 1813 2333 1836
rect 2338 1803 2341 1816
rect 2346 1813 2349 1843
rect 2378 1813 2381 2006
rect 2402 1996 2405 2053
rect 2434 2046 2437 2126
rect 2454 2106 2457 2163
rect 2418 2043 2437 2046
rect 2450 2103 2457 2106
rect 2418 2003 2421 2043
rect 2442 2023 2445 2036
rect 2450 2003 2453 2103
rect 2466 2036 2469 2156
rect 2490 2086 2493 2163
rect 2514 2103 2517 2126
rect 2462 2033 2469 2036
rect 2482 2083 2493 2086
rect 2538 2083 2541 2193
rect 2558 2156 2561 2263
rect 2666 2256 2669 2273
rect 2698 2266 2701 2326
rect 2738 2323 2749 2326
rect 2662 2253 2669 2256
rect 2674 2263 2709 2266
rect 2570 2176 2573 2216
rect 2610 2176 2613 2206
rect 2570 2173 2613 2176
rect 2558 2153 2565 2156
rect 2402 1993 2409 1996
rect 2406 1936 2409 1993
rect 2406 1933 2413 1936
rect 2418 1933 2421 1946
rect 2394 1893 2397 1916
rect 2410 1913 2413 1933
rect 2434 1846 2437 1996
rect 2462 1986 2465 2033
rect 2462 1983 2469 1986
rect 2466 1956 2469 1983
rect 2466 1953 2473 1956
rect 2458 1923 2461 1946
rect 2458 1886 2461 1916
rect 2454 1883 2461 1886
rect 2434 1843 2445 1846
rect 2434 1823 2437 1836
rect 2418 1813 2429 1816
rect 2346 1756 2349 1806
rect 2434 1796 2437 1806
rect 2330 1753 2349 1756
rect 2394 1793 2437 1796
rect 2306 1743 2317 1746
rect 2298 1733 2309 1736
rect 2298 1596 2301 1606
rect 2290 1593 2301 1596
rect 2250 1573 2261 1576
rect 2114 1423 2141 1426
rect 2114 1413 2133 1416
rect 2138 1406 2141 1423
rect 2130 1403 2141 1406
rect 2114 1213 2117 1336
rect 2130 1326 2133 1403
rect 2162 1376 2165 1406
rect 2178 1403 2181 1536
rect 2202 1523 2205 1573
rect 2226 1556 2229 1573
rect 2218 1553 2229 1556
rect 2218 1486 2221 1553
rect 2218 1483 2229 1486
rect 2226 1456 2229 1483
rect 2218 1453 2229 1456
rect 2250 1456 2253 1566
rect 2258 1553 2261 1573
rect 2290 1533 2293 1593
rect 2314 1546 2317 1743
rect 2330 1723 2333 1753
rect 2346 1686 2349 1736
rect 2394 1723 2397 1793
rect 2426 1723 2429 1736
rect 2442 1686 2445 1843
rect 2454 1766 2457 1883
rect 2470 1876 2473 1953
rect 2466 1873 2473 1876
rect 2454 1763 2461 1766
rect 2458 1693 2461 1763
rect 2346 1683 2445 1686
rect 2354 1576 2357 1646
rect 2370 1623 2373 1676
rect 2330 1573 2357 1576
rect 2386 1576 2389 1606
rect 2402 1603 2405 1683
rect 2466 1656 2469 1873
rect 2482 1836 2485 2083
rect 2562 2016 2565 2153
rect 2586 2103 2589 2126
rect 2602 2123 2613 2126
rect 2602 2036 2605 2123
rect 2610 2096 2613 2116
rect 2618 2103 2621 2236
rect 2634 2213 2645 2216
rect 2650 2206 2653 2216
rect 2634 2203 2653 2206
rect 2626 2163 2629 2196
rect 2626 2113 2629 2136
rect 2634 2133 2637 2203
rect 2662 2186 2665 2253
rect 2674 2203 2677 2263
rect 2698 2213 2701 2236
rect 2706 2213 2709 2263
rect 2662 2183 2669 2186
rect 2666 2163 2669 2183
rect 2722 2136 2725 2206
rect 2658 2096 2661 2126
rect 2706 2116 2709 2136
rect 2610 2093 2661 2096
rect 2698 2113 2709 2116
rect 2714 2133 2725 2136
rect 2738 2133 2741 2323
rect 2778 2303 2781 2373
rect 2802 2336 2805 2483
rect 2818 2436 2821 2666
rect 2826 2603 2829 2656
rect 2834 2603 2837 2723
rect 2858 2713 2861 2736
rect 2874 2723 2877 2763
rect 2890 2723 2893 2736
rect 2914 2723 2917 2746
rect 2970 2713 2973 2726
rect 2874 2613 2877 2626
rect 2898 2593 2901 2606
rect 2866 2563 2909 2566
rect 2866 2533 2869 2563
rect 2826 2493 2829 2526
rect 2882 2456 2885 2536
rect 2906 2523 2909 2563
rect 2954 2523 2965 2526
rect 2810 2433 2821 2436
rect 2874 2453 2885 2456
rect 2810 2366 2813 2433
rect 2850 2413 2853 2426
rect 2826 2393 2829 2406
rect 2874 2393 2877 2453
rect 2898 2413 2909 2416
rect 2946 2366 2949 2386
rect 2810 2363 2829 2366
rect 2802 2333 2813 2336
rect 2778 2216 2781 2226
rect 2754 2213 2765 2216
rect 2770 2213 2781 2216
rect 2754 2136 2757 2213
rect 2762 2136 2765 2146
rect 2754 2133 2765 2136
rect 2698 2036 2701 2113
rect 2602 2033 2653 2036
rect 2698 2033 2709 2036
rect 2530 1976 2533 2016
rect 2562 2013 2581 2016
rect 2586 2013 2597 2016
rect 2650 2013 2653 2033
rect 2554 2003 2573 2006
rect 2554 1976 2557 2003
rect 2530 1973 2557 1976
rect 2562 1993 2573 1996
rect 2562 1966 2565 1993
rect 2578 1976 2581 2013
rect 2626 1993 2629 2006
rect 2674 1983 2677 2006
rect 2546 1923 2549 1966
rect 2554 1963 2565 1966
rect 2554 1943 2557 1963
rect 2554 1896 2557 1936
rect 2562 1913 2565 1963
rect 2574 1973 2581 1976
rect 2574 1916 2577 1973
rect 2586 1923 2589 1966
rect 2574 1913 2581 1916
rect 2538 1893 2557 1896
rect 2482 1833 2493 1836
rect 2490 1776 2493 1833
rect 2538 1813 2541 1893
rect 2578 1826 2581 1913
rect 2570 1823 2581 1826
rect 2490 1773 2509 1776
rect 2474 1723 2477 1766
rect 2490 1733 2493 1746
rect 2506 1733 2509 1773
rect 2530 1723 2533 1746
rect 2466 1653 2473 1656
rect 2426 1576 2429 1616
rect 2386 1573 2429 1576
rect 2314 1543 2321 1546
rect 2274 1493 2277 1526
rect 2318 1496 2321 1543
rect 2314 1493 2321 1496
rect 2250 1453 2261 1456
rect 2202 1376 2205 1416
rect 2218 1406 2221 1453
rect 2218 1403 2229 1406
rect 2162 1373 2205 1376
rect 2146 1333 2165 1336
rect 2186 1333 2189 1356
rect 2122 1313 2125 1326
rect 2130 1323 2157 1326
rect 2162 1216 2165 1333
rect 2194 1306 2197 1346
rect 2210 1333 2213 1386
rect 2226 1346 2229 1403
rect 2258 1376 2261 1453
rect 2314 1436 2317 1493
rect 2330 1476 2333 1573
rect 2338 1563 2381 1566
rect 2338 1523 2341 1563
rect 2378 1533 2381 1563
rect 2386 1543 2389 1556
rect 2402 1523 2405 1546
rect 2458 1536 2461 1556
rect 2450 1533 2461 1536
rect 2330 1473 2341 1476
rect 2310 1433 2317 1436
rect 2290 1376 2293 1406
rect 2250 1373 2261 1376
rect 2282 1373 2293 1376
rect 2250 1356 2253 1373
rect 2246 1353 2253 1356
rect 2226 1343 2237 1346
rect 2194 1303 2205 1306
rect 2154 1213 2165 1216
rect 2186 1213 2197 1216
rect 2082 1146 2085 1173
rect 2154 1166 2157 1213
rect 2170 1183 2173 1206
rect 2154 1163 2165 1166
rect 2066 1123 2069 1146
rect 2078 1143 2085 1146
rect 2078 1086 2081 1143
rect 2130 1123 2133 1136
rect 2138 1103 2141 1136
rect 2146 1123 2149 1146
rect 2162 1106 2165 1163
rect 2202 1143 2205 1303
rect 2234 1243 2237 1343
rect 2246 1296 2249 1353
rect 2258 1323 2261 1336
rect 2246 1293 2253 1296
rect 2210 1213 2221 1216
rect 2210 1156 2213 1213
rect 2250 1196 2253 1293
rect 2282 1226 2285 1373
rect 2310 1366 2313 1433
rect 2322 1413 2325 1426
rect 2338 1376 2341 1473
rect 2298 1363 2313 1366
rect 2330 1373 2341 1376
rect 2298 1273 2301 1363
rect 2306 1353 2325 1356
rect 2306 1323 2309 1353
rect 2330 1343 2333 1373
rect 2282 1223 2293 1226
rect 2250 1193 2261 1196
rect 2290 1193 2293 1223
rect 2298 1213 2301 1236
rect 2306 1216 2309 1246
rect 2314 1226 2317 1336
rect 2330 1333 2341 1336
rect 2346 1333 2349 1356
rect 2378 1333 2381 1416
rect 2394 1373 2397 1406
rect 2426 1336 2429 1526
rect 2450 1466 2453 1533
rect 2470 1526 2473 1653
rect 2482 1613 2485 1656
rect 2514 1613 2525 1616
rect 2514 1596 2517 1613
rect 2466 1523 2473 1526
rect 2450 1463 2461 1466
rect 2418 1333 2429 1336
rect 2442 1333 2445 1416
rect 2458 1353 2461 1463
rect 2322 1306 2325 1326
rect 2322 1303 2329 1306
rect 2326 1236 2329 1303
rect 2326 1233 2333 1236
rect 2314 1223 2325 1226
rect 2306 1213 2317 1216
rect 2322 1213 2325 1223
rect 2330 1206 2333 1233
rect 2338 1216 2341 1266
rect 2346 1233 2349 1326
rect 2338 1213 2345 1216
rect 2306 1203 2333 1206
rect 2242 1166 2245 1186
rect 2242 1163 2249 1166
rect 2210 1153 2229 1156
rect 2210 1136 2213 1153
rect 2154 1103 2165 1106
rect 2078 1083 2085 1086
rect 2082 1016 2085 1083
rect 2074 1013 2085 1016
rect 2074 1003 2077 1013
rect 2106 993 2109 1006
rect 2122 1003 2125 1026
rect 2154 986 2157 1103
rect 2170 1013 2173 1136
rect 2178 1106 2181 1136
rect 2194 1133 2213 1136
rect 2218 1133 2221 1146
rect 2226 1133 2229 1153
rect 2194 1123 2197 1133
rect 2234 1126 2237 1136
rect 2202 1123 2213 1126
rect 2226 1123 2237 1126
rect 2202 1116 2205 1123
rect 2186 1113 2205 1116
rect 2226 1113 2229 1123
rect 2246 1116 2249 1163
rect 2242 1113 2249 1116
rect 2178 1103 2221 1106
rect 2210 1036 2213 1056
rect 2202 1033 2213 1036
rect 2154 983 2165 986
rect 2162 966 2165 983
rect 2074 963 2117 966
rect 2162 963 2173 966
rect 2074 933 2077 963
rect 2090 873 2093 936
rect 2114 923 2117 963
rect 2170 886 2173 963
rect 2162 883 2173 886
rect 2162 843 2165 883
rect 2202 846 2205 1033
rect 2218 853 2221 1103
rect 2226 1013 2229 1106
rect 2242 1053 2245 1113
rect 2258 1066 2261 1193
rect 2274 1136 2277 1176
rect 2306 1156 2309 1203
rect 2282 1153 2309 1156
rect 2282 1143 2285 1153
rect 2274 1133 2293 1136
rect 2290 1116 2293 1133
rect 2298 1123 2301 1146
rect 2306 1133 2309 1153
rect 2314 1123 2317 1156
rect 2290 1113 2301 1116
rect 2250 1063 2261 1066
rect 2250 1046 2253 1063
rect 2242 1043 2253 1046
rect 2226 913 2229 926
rect 2242 873 2245 1043
rect 2258 1003 2261 1026
rect 2290 1013 2293 1106
rect 2298 1073 2301 1113
rect 2202 843 2253 846
rect 2042 776 2045 816
rect 2002 773 2045 776
rect 1986 726 1989 736
rect 1978 723 1989 726
rect 2050 723 2053 746
rect 1978 716 1981 723
rect 1954 713 1981 716
rect 1930 703 1937 706
rect 1934 566 1937 703
rect 1954 666 1957 713
rect 1986 703 1989 716
rect 2058 706 2061 796
rect 2106 776 2109 816
rect 2106 773 2117 776
rect 2066 763 2109 766
rect 2066 733 2069 763
rect 2082 733 2085 746
rect 2106 723 2109 763
rect 2058 703 2077 706
rect 1946 663 1957 666
rect 1946 613 1949 663
rect 1978 613 1981 626
rect 2026 613 2037 616
rect 2050 606 2053 626
rect 1934 563 1965 566
rect 1914 553 1925 556
rect 1890 523 1893 546
rect 1882 513 1901 516
rect 1858 453 1877 456
rect 1858 396 1861 453
rect 1874 413 1877 436
rect 1834 333 1845 336
rect 1850 393 1861 396
rect 1850 326 1853 393
rect 1858 336 1861 376
rect 1890 346 1893 416
rect 1898 406 1901 513
rect 1906 413 1909 446
rect 1898 403 1909 406
rect 1882 343 1893 346
rect 1858 333 1877 336
rect 1786 313 1789 326
rect 1810 293 1813 326
rect 1730 213 1765 216
rect 1714 166 1717 183
rect 1706 163 1717 166
rect 1706 116 1709 163
rect 1730 123 1733 213
rect 1810 203 1813 216
rect 1818 213 1821 326
rect 1842 323 1853 326
rect 1842 266 1845 323
rect 1866 293 1869 326
rect 1834 263 1845 266
rect 1834 206 1837 263
rect 1874 246 1877 333
rect 1882 313 1885 343
rect 1874 243 1881 246
rect 1818 203 1837 206
rect 1746 133 1749 146
rect 1818 136 1821 203
rect 1850 193 1853 206
rect 1878 196 1881 243
rect 1890 213 1893 336
rect 1906 293 1909 403
rect 1914 333 1917 553
rect 1930 533 1933 556
rect 1962 456 1965 563
rect 1978 523 1981 556
rect 1930 453 1965 456
rect 2010 516 2013 526
rect 2018 523 2021 606
rect 2042 553 2045 606
rect 2050 603 2057 606
rect 2054 546 2057 603
rect 2050 543 2057 546
rect 2026 516 2029 536
rect 2010 513 2029 516
rect 1922 383 1925 406
rect 1930 376 1933 453
rect 1922 373 1933 376
rect 1922 326 1925 373
rect 1938 363 1941 416
rect 1954 413 1957 436
rect 2010 426 2013 513
rect 2050 486 2053 543
rect 2066 523 2069 616
rect 2074 583 2077 703
rect 2114 676 2117 773
rect 2122 743 2125 806
rect 2170 803 2173 816
rect 2170 753 2189 756
rect 2162 686 2165 726
rect 2106 673 2117 676
rect 2130 683 2165 686
rect 2106 556 2109 673
rect 2122 593 2125 616
rect 2130 586 2133 683
rect 2154 603 2157 676
rect 2170 603 2173 753
rect 2186 733 2189 753
rect 2210 686 2213 756
rect 2206 683 2213 686
rect 2130 583 2141 586
rect 2074 553 2109 556
rect 2042 483 2053 486
rect 2002 423 2037 426
rect 1914 323 1925 326
rect 1914 206 1917 323
rect 1922 293 1925 316
rect 1930 313 1933 326
rect 1946 313 1949 356
rect 1962 343 1965 416
rect 2002 403 2005 423
rect 2010 356 2013 416
rect 2026 403 2029 416
rect 1970 333 1973 356
rect 2010 353 2029 356
rect 1938 273 1941 306
rect 1994 293 1997 326
rect 2026 323 2029 353
rect 2034 333 2037 423
rect 2042 413 2045 436
rect 2074 416 2077 553
rect 2090 533 2093 546
rect 2106 513 2117 516
rect 2066 413 2077 416
rect 2042 326 2045 406
rect 2066 356 2069 413
rect 2090 373 2093 406
rect 2066 353 2077 356
rect 2058 333 2069 336
rect 2042 323 2053 326
rect 2058 306 2061 333
rect 2010 303 2061 306
rect 1922 213 1933 216
rect 2010 213 2013 303
rect 2034 216 2037 296
rect 2074 246 2077 353
rect 2082 306 2085 356
rect 2098 346 2101 416
rect 2090 343 2101 346
rect 2090 313 2093 343
rect 2106 323 2109 406
rect 2114 343 2117 416
rect 2122 373 2125 536
rect 2138 466 2141 583
rect 2162 516 2165 526
rect 2170 523 2173 546
rect 2194 543 2197 616
rect 2206 606 2209 683
rect 2202 603 2209 606
rect 2202 543 2205 603
rect 2218 556 2221 816
rect 2226 793 2229 806
rect 2234 783 2237 796
rect 2250 766 2253 843
rect 2258 813 2261 926
rect 2250 763 2257 766
rect 2226 673 2229 726
rect 2242 666 2245 686
rect 2238 663 2245 666
rect 2238 566 2241 663
rect 2254 656 2257 763
rect 2210 553 2221 556
rect 2234 563 2241 566
rect 2250 653 2257 656
rect 2162 513 2173 516
rect 2130 463 2141 466
rect 2122 336 2125 356
rect 2114 333 2125 336
rect 2130 336 2133 463
rect 2170 413 2173 513
rect 2210 456 2213 553
rect 2218 523 2221 546
rect 2210 453 2217 456
rect 2146 353 2149 406
rect 2130 333 2141 336
rect 2082 303 2101 306
rect 2066 243 2077 246
rect 2034 213 2045 216
rect 1914 203 1925 206
rect 1874 193 1881 196
rect 1842 143 1845 156
rect 1814 133 1821 136
rect 1706 113 1717 116
rect 1666 103 1677 106
rect 1650 83 1657 86
rect 1626 73 1637 76
rect 1634 0 1637 73
rect 1650 0 1653 83
rect 1666 0 1669 16
rect 1674 3 1677 103
rect 1674 0 1685 3
rect 1714 0 1717 113
rect 1746 0 1749 126
rect 1794 113 1797 126
rect 1814 76 1817 133
rect 1810 73 1817 76
rect 1826 76 1829 126
rect 1842 113 1845 136
rect 1874 123 1877 193
rect 1922 146 1925 203
rect 1962 193 1965 206
rect 1946 163 1989 166
rect 1898 133 1901 146
rect 1922 143 1933 146
rect 1930 96 1933 143
rect 1946 123 1949 163
rect 1986 133 1989 163
rect 2018 143 2021 156
rect 2042 146 2045 213
rect 2066 196 2069 243
rect 2082 213 2085 236
rect 2090 203 2093 226
rect 2066 193 2077 196
rect 2034 143 2045 146
rect 2066 143 2069 156
rect 1914 93 1933 96
rect 1826 73 1837 76
rect 1810 16 1813 73
rect 1810 13 1821 16
rect 1818 0 1821 13
rect 1834 0 1837 73
rect 1914 0 1917 93
rect 1978 0 1981 126
rect 2034 123 2037 143
rect 2074 116 2077 193
rect 2098 123 2101 303
rect 2114 193 2117 333
rect 2122 313 2125 326
rect 2130 233 2133 326
rect 2138 253 2141 333
rect 2146 316 2149 336
rect 2202 333 2205 376
rect 2214 356 2217 453
rect 2234 436 2237 563
rect 2234 433 2245 436
rect 2226 373 2229 416
rect 2242 403 2245 433
rect 2250 383 2253 653
rect 2266 613 2269 846
rect 2282 796 2285 1006
rect 2298 996 2301 1066
rect 2294 993 2301 996
rect 2294 906 2297 993
rect 2306 976 2309 1026
rect 2322 1003 2325 1196
rect 2330 1133 2333 1166
rect 2342 1086 2345 1213
rect 2354 1153 2357 1276
rect 2362 1213 2365 1326
rect 2370 1313 2373 1326
rect 2442 1253 2445 1316
rect 2458 1243 2461 1346
rect 2466 1333 2469 1523
rect 2482 1496 2485 1596
rect 2490 1553 2493 1596
rect 2506 1593 2517 1596
rect 2506 1536 2509 1593
rect 2522 1576 2525 1606
rect 2538 1603 2541 1656
rect 2570 1626 2573 1823
rect 2578 1803 2581 1816
rect 2594 1776 2597 1806
rect 2626 1776 2629 1976
rect 2682 1966 2685 2006
rect 2690 2003 2693 2016
rect 2698 1966 2701 1986
rect 2658 1963 2685 1966
rect 2694 1963 2701 1966
rect 2658 1916 2661 1963
rect 2674 1923 2677 1956
rect 2658 1913 2669 1916
rect 2642 1783 2645 1816
rect 2666 1793 2669 1913
rect 2694 1876 2697 1963
rect 2706 1923 2709 2033
rect 2714 1966 2717 2133
rect 2722 2013 2725 2126
rect 2730 2123 2741 2126
rect 2730 2113 2733 2123
rect 2754 2083 2757 2126
rect 2762 2106 2765 2133
rect 2770 2113 2773 2213
rect 2786 2203 2789 2216
rect 2802 2203 2805 2326
rect 2810 2316 2813 2333
rect 2810 2313 2817 2316
rect 2814 2196 2817 2313
rect 2826 2286 2829 2363
rect 2858 2323 2861 2366
rect 2938 2363 2949 2366
rect 2826 2283 2837 2286
rect 2810 2193 2817 2196
rect 2826 2193 2829 2206
rect 2762 2103 2773 2106
rect 2762 2013 2765 2036
rect 2770 2006 2773 2103
rect 2778 2013 2781 2136
rect 2786 2093 2789 2126
rect 2722 1983 2725 2006
rect 2762 2003 2773 2006
rect 2794 1996 2797 2136
rect 2770 1993 2797 1996
rect 2802 1993 2805 2006
rect 2714 1963 2721 1966
rect 2718 1916 2721 1963
rect 2730 1933 2733 1946
rect 2754 1933 2757 1956
rect 2690 1873 2697 1876
rect 2714 1913 2721 1916
rect 2594 1773 2629 1776
rect 2690 1776 2693 1873
rect 2714 1836 2717 1913
rect 2738 1846 2741 1926
rect 2762 1923 2765 1946
rect 2770 1933 2773 1993
rect 2810 1926 2813 2193
rect 2826 2133 2829 2146
rect 2818 2113 2821 2126
rect 2834 2106 2837 2283
rect 2842 2133 2845 2216
rect 2866 2203 2869 2306
rect 2938 2266 2941 2363
rect 2938 2263 2945 2266
rect 2858 2123 2861 2146
rect 2898 2136 2901 2216
rect 2942 2166 2945 2263
rect 2954 2193 2957 2216
rect 2938 2163 2945 2166
rect 2898 2133 2909 2136
rect 2898 2113 2909 2116
rect 2826 2103 2837 2106
rect 2826 1946 2829 2103
rect 2938 2066 2941 2163
rect 2938 2063 2949 2066
rect 2946 2046 2949 2063
rect 2866 2023 2869 2036
rect 2858 2013 2869 2016
rect 2858 2006 2861 2013
rect 2842 2003 2861 2006
rect 2866 1993 2869 2006
rect 2874 2003 2877 2046
rect 2946 2043 2953 2046
rect 2914 1973 2917 2006
rect 2938 1993 2941 2016
rect 2802 1923 2813 1926
rect 2818 1943 2829 1946
rect 2866 1963 2909 1966
rect 2754 1856 2757 1916
rect 2754 1853 2761 1856
rect 2738 1843 2749 1846
rect 2706 1833 2741 1836
rect 2706 1813 2709 1833
rect 2722 1823 2733 1826
rect 2706 1793 2709 1806
rect 2714 1776 2717 1816
rect 2722 1813 2733 1816
rect 2722 1793 2725 1813
rect 2730 1783 2733 1806
rect 2738 1803 2741 1833
rect 2746 1776 2749 1843
rect 2758 1776 2761 1853
rect 2690 1773 2701 1776
rect 2594 1683 2597 1726
rect 2610 1723 2613 1773
rect 2658 1723 2661 1746
rect 2570 1623 2581 1626
rect 2562 1576 2565 1616
rect 2522 1573 2565 1576
rect 2490 1533 2509 1536
rect 2506 1526 2509 1533
rect 2498 1503 2501 1526
rect 2506 1523 2517 1526
rect 2506 1513 2517 1516
rect 2506 1496 2509 1513
rect 2482 1493 2509 1496
rect 2474 1393 2477 1416
rect 2482 1263 2485 1493
rect 2522 1413 2525 1536
rect 2546 1456 2549 1536
rect 2562 1503 2565 1526
rect 2578 1496 2581 1623
rect 2634 1603 2637 1616
rect 2642 1603 2645 1646
rect 2610 1533 2637 1536
rect 2634 1523 2637 1533
rect 2570 1493 2581 1496
rect 2570 1473 2573 1493
rect 2546 1453 2581 1456
rect 2546 1436 2549 1453
rect 2538 1433 2549 1436
rect 2498 1373 2501 1406
rect 2538 1366 2541 1433
rect 2578 1413 2581 1453
rect 2642 1413 2645 1536
rect 2650 1503 2653 1616
rect 2658 1453 2661 1676
rect 2666 1563 2669 1626
rect 2674 1576 2677 1606
rect 2690 1603 2693 1726
rect 2698 1723 2701 1773
rect 2714 1773 2749 1776
rect 2754 1773 2761 1776
rect 2714 1663 2717 1773
rect 2722 1733 2741 1736
rect 2746 1733 2749 1746
rect 2738 1726 2741 1733
rect 2738 1723 2749 1726
rect 2738 1713 2749 1716
rect 2722 1686 2725 1706
rect 2722 1683 2733 1686
rect 2714 1576 2717 1616
rect 2674 1573 2717 1576
rect 2730 1566 2733 1683
rect 2754 1566 2757 1773
rect 2770 1766 2773 1856
rect 2802 1826 2805 1923
rect 2818 1906 2821 1943
rect 2866 1933 2869 1963
rect 2826 1923 2845 1926
rect 2818 1903 2829 1906
rect 2826 1846 2829 1903
rect 2882 1856 2885 1956
rect 2906 1923 2909 1963
rect 2950 1946 2953 2043
rect 2946 1943 2953 1946
rect 2794 1823 2805 1826
rect 2818 1843 2829 1846
rect 2874 1853 2885 1856
rect 2818 1823 2821 1843
rect 2794 1796 2797 1823
rect 2810 1813 2829 1816
rect 2858 1803 2861 1826
rect 2794 1793 2805 1796
rect 2770 1763 2777 1766
rect 2762 1733 2765 1756
rect 2774 1706 2777 1763
rect 2770 1703 2777 1706
rect 2786 1703 2789 1786
rect 2770 1686 2773 1703
rect 2802 1696 2805 1793
rect 2858 1733 2861 1746
rect 2874 1733 2877 1853
rect 2898 1813 2901 1826
rect 2818 1723 2837 1726
rect 2898 1723 2901 1746
rect 2714 1563 2733 1566
rect 2746 1563 2757 1566
rect 2762 1683 2773 1686
rect 2798 1693 2805 1696
rect 2714 1543 2717 1563
rect 2674 1533 2693 1536
rect 2690 1413 2693 1533
rect 2714 1523 2733 1526
rect 2746 1516 2749 1563
rect 2730 1513 2749 1516
rect 2730 1426 2733 1513
rect 2762 1496 2765 1683
rect 2770 1606 2773 1616
rect 2778 1613 2781 1636
rect 2770 1603 2781 1606
rect 2770 1506 2773 1536
rect 2786 1533 2789 1646
rect 2798 1626 2801 1693
rect 2946 1656 2949 1943
rect 2962 1936 2965 2396
rect 2986 2186 2989 2446
rect 2986 2183 2997 2186
rect 2978 1953 2981 2176
rect 2994 2066 2997 2183
rect 2986 2063 2997 2066
rect 2986 1996 2989 2063
rect 2994 2013 2997 2046
rect 2986 1993 2997 1996
rect 2962 1933 2973 1936
rect 2954 1923 2965 1926
rect 2970 1886 2973 1933
rect 2962 1883 2973 1886
rect 2954 1723 2957 1736
rect 2946 1653 2953 1656
rect 2794 1623 2801 1626
rect 2794 1573 2797 1623
rect 2818 1613 2837 1616
rect 2802 1603 2829 1606
rect 2818 1573 2821 1596
rect 2770 1503 2781 1506
rect 2810 1503 2813 1526
rect 2762 1493 2773 1496
rect 2722 1423 2733 1426
rect 2610 1373 2613 1406
rect 2722 1366 2725 1423
rect 2538 1363 2549 1366
rect 2410 1193 2413 1206
rect 2426 1193 2429 1226
rect 2442 1223 2445 1236
rect 2362 1113 2365 1146
rect 2378 1113 2381 1136
rect 2362 1103 2373 1106
rect 2410 1093 2413 1126
rect 2342 1083 2349 1086
rect 2346 996 2349 1083
rect 2426 1043 2429 1136
rect 2434 1016 2437 1166
rect 2482 1133 2485 1176
rect 2498 1153 2501 1356
rect 2514 1256 2517 1346
rect 2546 1333 2549 1363
rect 2554 1336 2557 1366
rect 2722 1363 2733 1366
rect 2626 1343 2661 1346
rect 2554 1333 2573 1336
rect 2626 1333 2629 1343
rect 2658 1336 2661 1343
rect 2538 1313 2541 1326
rect 2510 1253 2517 1256
rect 2510 1196 2513 1253
rect 2522 1213 2525 1246
rect 2546 1243 2549 1326
rect 2510 1193 2517 1196
rect 2514 1173 2517 1193
rect 2418 1013 2437 1016
rect 2442 1006 2445 1076
rect 2466 1073 2469 1126
rect 2498 1106 2501 1146
rect 2522 1123 2525 1206
rect 2530 1183 2533 1206
rect 2538 1166 2541 1226
rect 2554 1213 2557 1333
rect 2650 1326 2653 1336
rect 2658 1333 2669 1336
rect 2722 1333 2725 1346
rect 2562 1303 2565 1326
rect 2570 1213 2573 1246
rect 2534 1163 2541 1166
rect 2482 1103 2501 1106
rect 2338 993 2349 996
rect 2306 973 2317 976
rect 2294 903 2301 906
rect 2274 793 2285 796
rect 2274 683 2277 793
rect 2282 743 2285 786
rect 2298 726 2301 903
rect 2314 833 2317 973
rect 2338 946 2341 993
rect 2402 976 2405 996
rect 2394 973 2405 976
rect 2338 943 2349 946
rect 2346 896 2349 943
rect 2362 923 2365 946
rect 2338 893 2349 896
rect 2330 813 2333 826
rect 2306 803 2317 806
rect 2330 733 2333 746
rect 2290 723 2301 726
rect 2290 636 2293 723
rect 2290 633 2301 636
rect 2258 486 2261 606
rect 2274 533 2277 546
rect 2290 543 2293 616
rect 2298 496 2301 633
rect 2306 596 2309 726
rect 2322 626 2325 726
rect 2314 623 2325 626
rect 2338 623 2341 893
rect 2354 803 2357 836
rect 2378 803 2381 816
rect 2354 733 2357 796
rect 2378 723 2381 746
rect 2394 686 2397 973
rect 2418 783 2421 1006
rect 2434 1003 2445 1006
rect 2434 956 2437 1003
rect 2466 976 2469 1006
rect 2482 993 2485 1103
rect 2534 1096 2537 1163
rect 2534 1093 2541 1096
rect 2546 1093 2549 1196
rect 2538 1073 2541 1093
rect 2570 1086 2573 1156
rect 2578 1133 2581 1326
rect 2642 1323 2653 1326
rect 2642 1213 2645 1323
rect 2650 1303 2653 1316
rect 2666 1216 2669 1333
rect 2730 1253 2733 1363
rect 2666 1213 2693 1216
rect 2698 1213 2701 1246
rect 2738 1213 2741 1416
rect 2754 1413 2757 1446
rect 2770 1413 2773 1493
rect 2746 1363 2749 1406
rect 2754 1323 2765 1326
rect 2754 1293 2757 1316
rect 2762 1313 2773 1316
rect 2778 1286 2781 1406
rect 2826 1396 2829 1603
rect 2866 1576 2869 1606
rect 2882 1603 2885 1646
rect 2906 1576 2909 1616
rect 2950 1576 2953 1653
rect 2962 1643 2965 1883
rect 2994 1876 2997 1993
rect 2986 1873 2997 1876
rect 2962 1613 2965 1636
rect 2866 1573 2909 1576
rect 2946 1573 2953 1576
rect 2986 1576 2989 1873
rect 3010 1813 3013 1826
rect 2986 1573 2997 1576
rect 2946 1456 2949 1573
rect 2978 1533 2981 1566
rect 2994 1526 2997 1573
rect 2986 1523 2997 1526
rect 2942 1453 2949 1456
rect 2858 1423 2861 1446
rect 2834 1403 2853 1406
rect 2826 1393 2845 1396
rect 2794 1296 2797 1336
rect 2818 1313 2821 1326
rect 2794 1293 2805 1296
rect 2762 1283 2781 1286
rect 2594 1166 2597 1206
rect 2690 1186 2693 1213
rect 2746 1203 2749 1276
rect 2754 1213 2757 1246
rect 2762 1203 2765 1283
rect 2770 1213 2773 1266
rect 2778 1206 2781 1256
rect 2802 1226 2805 1293
rect 2842 1273 2845 1393
rect 2850 1286 2853 1403
rect 2882 1376 2885 1406
rect 2898 1393 2901 1406
rect 2922 1376 2925 1416
rect 2882 1373 2925 1376
rect 2898 1333 2901 1366
rect 2922 1333 2925 1366
rect 2930 1326 2933 1396
rect 2942 1376 2945 1453
rect 2962 1436 2965 1456
rect 2962 1433 2969 1436
rect 2966 1376 2969 1433
rect 2986 1426 2989 1523
rect 3010 1483 3013 1526
rect 2986 1423 2997 1426
rect 2942 1373 2949 1376
rect 2874 1293 2877 1326
rect 2882 1286 2885 1326
rect 2922 1323 2933 1326
rect 2850 1283 2893 1286
rect 2770 1203 2781 1206
rect 2794 1223 2805 1226
rect 2850 1223 2853 1246
rect 2794 1203 2797 1223
rect 2826 1213 2853 1216
rect 2826 1203 2829 1213
rect 2690 1183 2701 1186
rect 2594 1163 2621 1166
rect 2594 1133 2597 1146
rect 2578 1103 2581 1126
rect 2570 1083 2581 1086
rect 2506 976 2509 1016
rect 2570 993 2573 1016
rect 2578 993 2581 1083
rect 2594 1013 2597 1116
rect 2618 1043 2621 1163
rect 2626 1126 2629 1166
rect 2642 1163 2693 1166
rect 2626 1123 2633 1126
rect 2642 1123 2645 1163
rect 2630 1066 2633 1123
rect 2626 1063 2633 1066
rect 2466 973 2509 976
rect 2610 976 2613 1006
rect 2626 1003 2629 1063
rect 2650 976 2653 1016
rect 2610 973 2653 976
rect 2658 966 2661 1136
rect 2674 1123 2677 1146
rect 2682 1143 2685 1156
rect 2690 1133 2693 1163
rect 2698 1123 2701 1183
rect 2730 1133 2733 1166
rect 2754 1156 2757 1176
rect 2754 1153 2761 1156
rect 2758 1096 2761 1153
rect 2754 1093 2761 1096
rect 2650 963 2661 966
rect 2650 956 2653 963
rect 2434 953 2477 956
rect 2434 923 2437 953
rect 2442 933 2461 936
rect 2466 933 2469 946
rect 2474 933 2477 953
rect 2618 953 2653 956
rect 2458 926 2461 933
rect 2426 816 2429 856
rect 2426 813 2437 816
rect 2426 723 2437 726
rect 2394 683 2413 686
rect 2314 613 2317 623
rect 2410 616 2413 683
rect 2442 623 2445 856
rect 2450 816 2453 926
rect 2458 923 2485 926
rect 2466 903 2469 916
rect 2482 896 2485 923
rect 2618 906 2621 953
rect 2650 933 2653 946
rect 2618 903 2629 906
rect 2482 893 2509 896
rect 2450 813 2461 816
rect 2458 723 2461 813
rect 2466 783 2469 796
rect 2474 733 2477 746
rect 2490 716 2493 876
rect 2506 836 2509 893
rect 2498 833 2509 836
rect 2498 813 2501 833
rect 2506 743 2509 786
rect 2530 776 2533 806
rect 2546 793 2549 806
rect 2570 776 2573 816
rect 2530 773 2573 776
rect 2626 766 2629 903
rect 2666 826 2669 836
rect 2674 826 2677 1046
rect 2738 1013 2741 1026
rect 2698 923 2701 966
rect 2738 956 2741 1006
rect 2746 996 2749 1016
rect 2754 996 2757 1093
rect 2770 1023 2773 1203
rect 2778 1163 2797 1166
rect 2778 1123 2781 1163
rect 2794 1136 2797 1163
rect 2826 1136 2829 1166
rect 2834 1146 2837 1156
rect 2834 1143 2845 1146
rect 2794 1133 2821 1136
rect 2826 1133 2837 1136
rect 2826 1083 2829 1126
rect 2746 993 2757 996
rect 2738 953 2749 956
rect 2738 906 2741 926
rect 2746 923 2749 953
rect 2730 903 2741 906
rect 2666 823 2677 826
rect 2682 833 2709 836
rect 2562 763 2605 766
rect 2490 713 2501 716
rect 2322 613 2341 616
rect 2410 613 2417 616
rect 2506 613 2509 736
rect 2538 646 2541 746
rect 2562 733 2565 763
rect 2538 643 2549 646
rect 2322 603 2341 606
rect 2306 593 2313 596
rect 2310 506 2313 593
rect 2322 523 2325 603
rect 2310 503 2317 506
rect 2290 493 2301 496
rect 2258 483 2269 486
rect 2266 436 2269 483
rect 2258 433 2269 436
rect 2258 406 2261 433
rect 2266 413 2277 416
rect 2258 403 2269 406
rect 2210 353 2217 356
rect 2210 326 2213 353
rect 2146 313 2157 316
rect 2154 213 2157 313
rect 2186 293 2189 326
rect 2202 323 2213 326
rect 2162 236 2165 256
rect 2162 233 2173 236
rect 2130 193 2133 206
rect 2114 163 2157 166
rect 2114 133 2117 163
rect 2130 133 2133 146
rect 2154 123 2157 163
rect 2170 116 2173 233
rect 2074 113 2101 116
rect 2098 0 2101 113
rect 2162 113 2173 116
rect 2162 0 2165 113
rect 2202 76 2205 323
rect 2218 256 2221 336
rect 2266 333 2269 403
rect 2218 253 2229 256
rect 2210 213 2213 226
rect 2226 173 2229 253
rect 2234 203 2237 226
rect 2250 186 2253 326
rect 2266 273 2269 326
rect 2274 313 2277 336
rect 2282 316 2285 416
rect 2290 406 2293 493
rect 2298 413 2301 456
rect 2314 426 2317 503
rect 2338 476 2341 546
rect 2306 423 2317 426
rect 2330 473 2341 476
rect 2290 403 2301 406
rect 2298 323 2301 403
rect 2306 323 2309 423
rect 2314 383 2317 406
rect 2330 356 2333 473
rect 2346 366 2349 576
rect 2386 533 2389 546
rect 2402 543 2405 606
rect 2354 503 2357 526
rect 2414 476 2417 613
rect 2538 606 2541 616
rect 2546 613 2549 643
rect 2578 636 2581 756
rect 2602 723 2605 763
rect 2618 763 2629 766
rect 2618 686 2621 763
rect 2618 683 2629 686
rect 2578 633 2589 636
rect 2426 523 2429 606
rect 2458 553 2461 606
rect 2538 603 2549 606
rect 2586 603 2589 633
rect 2414 473 2429 476
rect 2370 423 2405 426
rect 2370 416 2373 423
rect 2354 393 2357 416
rect 2362 413 2373 416
rect 2386 403 2389 416
rect 2402 413 2405 423
rect 2378 393 2397 396
rect 2346 363 2357 366
rect 2330 353 2341 356
rect 2282 313 2317 316
rect 2322 296 2325 336
rect 2314 293 2325 296
rect 2314 213 2317 293
rect 2338 256 2341 353
rect 2334 253 2341 256
rect 2266 193 2269 206
rect 2334 186 2337 253
rect 2354 246 2357 363
rect 2370 323 2381 326
rect 2370 293 2373 323
rect 2378 313 2389 316
rect 2394 313 2397 393
rect 2426 366 2429 473
rect 2450 403 2453 436
rect 2466 406 2469 526
rect 2506 523 2509 546
rect 2458 403 2469 406
rect 2410 363 2429 366
rect 2386 293 2389 306
rect 2346 243 2357 246
rect 2250 183 2261 186
rect 2334 183 2341 186
rect 2218 143 2221 156
rect 2194 73 2205 76
rect 2194 16 2197 73
rect 2194 13 2205 16
rect 2202 0 2205 13
rect 2218 0 2221 126
rect 2258 116 2261 183
rect 2274 123 2277 176
rect 2290 163 2333 166
rect 2290 133 2293 163
rect 2306 133 2309 146
rect 2330 123 2333 163
rect 2258 113 2269 116
rect 2266 86 2269 113
rect 2266 83 2277 86
rect 2250 0 2253 76
rect 2274 16 2277 83
rect 2338 73 2341 183
rect 2346 153 2349 243
rect 2402 233 2405 336
rect 2410 296 2413 363
rect 2458 333 2461 403
rect 2434 313 2437 326
rect 2442 306 2445 326
rect 2474 316 2477 416
rect 2482 396 2485 406
rect 2490 403 2493 466
rect 2498 413 2501 426
rect 2482 393 2493 396
rect 2538 393 2541 603
rect 2554 543 2557 566
rect 2610 546 2613 616
rect 2626 566 2629 683
rect 2650 626 2653 806
rect 2666 786 2669 823
rect 2674 793 2677 816
rect 2682 813 2685 833
rect 2698 813 2701 826
rect 2706 813 2709 833
rect 2666 783 2677 786
rect 2674 733 2677 783
rect 2658 703 2661 726
rect 2698 723 2701 806
rect 2730 796 2733 903
rect 2746 803 2749 826
rect 2754 813 2757 993
rect 2762 963 2765 1006
rect 2834 1003 2837 1133
rect 2842 1116 2845 1143
rect 2850 1123 2853 1213
rect 2858 1203 2861 1236
rect 2890 1226 2893 1283
rect 2922 1276 2925 1323
rect 2914 1273 2925 1276
rect 2890 1223 2901 1226
rect 2874 1193 2877 1206
rect 2858 1116 2861 1146
rect 2842 1113 2861 1116
rect 2882 1013 2885 1126
rect 2898 1123 2901 1223
rect 2914 1126 2917 1273
rect 2938 1213 2941 1236
rect 2914 1123 2925 1126
rect 2922 966 2925 1123
rect 2946 1033 2949 1373
rect 2962 1373 2969 1376
rect 2962 1256 2965 1373
rect 2978 1363 2981 1416
rect 2994 1356 2997 1423
rect 2986 1353 2997 1356
rect 2986 1276 2989 1353
rect 2958 1253 2965 1256
rect 2982 1273 2989 1276
rect 2958 1176 2961 1253
rect 2982 1186 2985 1273
rect 2994 1263 3005 1266
rect 3002 1246 3005 1263
rect 3002 1243 3009 1246
rect 2994 1193 2997 1216
rect 3006 1186 3009 1243
rect 2982 1183 2989 1186
rect 2958 1173 2965 1176
rect 2842 963 2885 966
rect 2922 963 2929 966
rect 2786 906 2789 946
rect 2842 933 2845 963
rect 2794 923 2813 926
rect 2730 793 2741 796
rect 2650 623 2677 626
rect 2738 623 2741 793
rect 2770 773 2773 906
rect 2786 903 2797 906
rect 2794 826 2797 903
rect 2858 876 2861 936
rect 2882 923 2885 963
rect 2926 906 2929 963
rect 2922 903 2929 906
rect 2938 903 2941 926
rect 2922 886 2925 903
rect 2906 883 2925 886
rect 2858 873 2869 876
rect 2786 823 2797 826
rect 2786 793 2789 823
rect 2770 733 2773 746
rect 2746 723 2757 726
rect 2794 723 2797 806
rect 2818 766 2821 796
rect 2810 763 2821 766
rect 2658 613 2669 616
rect 2674 613 2677 623
rect 2722 613 2741 616
rect 2746 606 2749 723
rect 2810 686 2813 763
rect 2834 756 2837 826
rect 2850 776 2853 806
rect 2866 803 2869 873
rect 2890 776 2893 816
rect 2850 773 2893 776
rect 2906 776 2909 883
rect 2962 853 2965 1173
rect 2986 836 2989 1183
rect 2978 833 2989 836
rect 3002 1183 3009 1186
rect 2938 813 2949 816
rect 2906 773 2917 776
rect 2834 753 2861 756
rect 2850 716 2853 726
rect 2858 723 2861 753
rect 2866 716 2869 736
rect 2850 713 2869 716
rect 2810 683 2821 686
rect 2706 603 2749 606
rect 2626 563 2637 566
rect 2570 523 2573 546
rect 2602 543 2613 546
rect 2610 516 2613 536
rect 2618 523 2621 536
rect 2602 513 2613 516
rect 2602 456 2605 513
rect 2634 506 2637 563
rect 2706 546 2709 603
rect 2722 563 2725 596
rect 2658 533 2661 546
rect 2706 543 2717 546
rect 2658 513 2661 526
rect 2682 506 2685 526
rect 2690 513 2693 526
rect 2626 503 2637 506
rect 2658 503 2685 506
rect 2602 453 2613 456
rect 2626 453 2629 503
rect 2610 436 2613 453
rect 2594 433 2613 436
rect 2490 326 2493 393
rect 2490 323 2517 326
rect 2474 313 2517 316
rect 2426 303 2445 306
rect 2410 293 2417 296
rect 2354 213 2357 226
rect 2402 203 2405 226
rect 2414 196 2417 293
rect 2410 193 2417 196
rect 2394 143 2397 156
rect 2410 143 2413 193
rect 2426 176 2429 303
rect 2522 256 2525 336
rect 2546 316 2549 416
rect 2562 323 2565 406
rect 2570 346 2573 406
rect 2586 353 2589 426
rect 2594 383 2597 433
rect 2658 423 2661 503
rect 2642 393 2645 406
rect 2666 403 2669 436
rect 2674 423 2677 436
rect 2714 433 2717 543
rect 2722 506 2725 526
rect 2722 503 2733 506
rect 2730 456 2733 503
rect 2722 453 2733 456
rect 2722 413 2725 453
rect 2730 413 2741 416
rect 2570 343 2629 346
rect 2570 333 2573 343
rect 2546 313 2597 316
rect 2602 296 2605 336
rect 2490 253 2525 256
rect 2586 293 2605 296
rect 2490 213 2493 253
rect 2522 213 2525 226
rect 2586 213 2589 293
rect 2626 236 2629 343
rect 2642 256 2645 336
rect 2698 333 2701 406
rect 2666 293 2669 326
rect 2642 253 2653 256
rect 2626 233 2637 236
rect 2634 216 2637 233
rect 2602 213 2637 216
rect 2650 213 2653 253
rect 2442 193 2445 206
rect 2538 193 2541 206
rect 2426 173 2445 176
rect 2266 13 2277 16
rect 2266 0 2269 13
rect 2386 0 2389 126
rect 2442 123 2445 173
rect 2466 163 2509 166
rect 2466 133 2469 163
rect 2482 133 2485 146
rect 2506 123 2509 163
rect 2570 143 2573 156
rect 2562 0 2565 126
rect 2602 123 2605 213
rect 2690 203 2693 226
rect 2610 163 2653 166
rect 2610 133 2613 163
rect 2626 133 2629 146
rect 2650 123 2653 163
rect 2706 156 2709 336
rect 2730 316 2733 413
rect 2746 326 2749 536
rect 2754 533 2757 626
rect 2770 576 2773 606
rect 2786 603 2789 636
rect 2810 576 2813 616
rect 2770 573 2813 576
rect 2818 563 2821 683
rect 2850 656 2853 713
rect 2850 653 2861 656
rect 2858 576 2861 653
rect 2850 573 2861 576
rect 2850 556 2853 573
rect 2842 553 2853 556
rect 2762 533 2773 536
rect 2778 533 2781 546
rect 2818 533 2829 536
rect 2762 503 2765 526
rect 2778 463 2781 526
rect 2754 413 2757 456
rect 2762 413 2765 436
rect 2810 383 2813 406
rect 2746 323 2765 326
rect 2730 313 2765 316
rect 2770 213 2773 336
rect 2818 316 2821 416
rect 2826 403 2829 533
rect 2842 496 2845 553
rect 2858 526 2861 536
rect 2866 533 2869 546
rect 2858 523 2869 526
rect 2874 523 2877 536
rect 2858 503 2861 516
rect 2842 493 2853 496
rect 2834 413 2837 426
rect 2834 336 2837 406
rect 2850 383 2853 493
rect 2866 356 2869 523
rect 2914 476 2917 773
rect 2938 523 2941 546
rect 2954 476 2957 776
rect 2978 736 2981 833
rect 2978 733 2989 736
rect 2986 713 2989 733
rect 2986 593 2989 616
rect 2986 523 2997 526
rect 2914 473 2941 476
rect 2954 473 2965 476
rect 2922 383 2925 406
rect 2930 403 2933 416
rect 2938 376 2941 473
rect 2962 376 2965 473
rect 3002 426 3005 1183
rect 3010 1013 3013 1036
rect 2994 423 3005 426
rect 2858 353 2869 356
rect 2914 373 2941 376
rect 2954 373 2965 376
rect 2826 333 2853 336
rect 2850 323 2853 333
rect 2858 326 2861 353
rect 2866 333 2869 346
rect 2858 323 2869 326
rect 2818 313 2853 316
rect 2866 296 2869 323
rect 2874 313 2877 336
rect 2858 293 2869 296
rect 2858 236 2861 293
rect 2858 233 2869 236
rect 2802 213 2805 226
rect 2866 213 2869 233
rect 2722 193 2725 206
rect 2882 196 2885 326
rect 2914 213 2917 373
rect 2938 323 2941 346
rect 2746 163 2789 166
rect 2706 153 2725 156
rect 2722 126 2725 153
rect 2730 143 2733 156
rect 2746 133 2749 163
rect 2762 133 2765 146
rect 2706 0 2709 126
rect 2722 123 2749 126
rect 2786 123 2789 163
rect 2850 156 2853 196
rect 2842 153 2853 156
rect 2850 143 2853 153
rect 2874 193 2885 196
rect 2898 193 2901 206
rect 2874 146 2877 193
rect 2874 143 2885 146
rect 2842 0 2845 126
rect 2882 123 2885 143
rect 2898 133 2901 146
rect 2914 133 2917 206
rect 2938 193 2941 216
rect 2938 123 2941 146
rect 2954 23 2957 373
rect 2994 313 2997 326
rect 2986 213 2997 216
rect 2986 123 2997 126
rect 3022 37 3042 3003
rect 3034 6 3037 26
rect 3046 13 3066 3027
rect 3074 6 3077 1716
rect 3034 3 3077 6
<< metal3 >>
rect 113 3032 1318 3037
rect 113 3022 118 3032
rect 1313 3027 1318 3032
rect 1313 3022 1526 3027
rect 41 3012 102 3017
rect 97 3007 102 3012
rect 329 3012 542 3017
rect 329 3007 334 3012
rect 97 3002 334 3007
rect 1473 3002 1566 3007
rect 353 2992 382 2997
rect 377 2987 382 2992
rect 553 2992 1454 2997
rect 553 2987 558 2992
rect 377 2982 558 2987
rect 1473 2977 1478 3002
rect 1561 2997 1566 3002
rect 1561 2992 1750 2997
rect 1497 2982 1550 2987
rect 1689 2982 1742 2987
rect 1313 2972 1478 2977
rect 1521 2972 1590 2977
rect 2097 2972 2206 2977
rect 761 2962 862 2967
rect 761 2957 766 2962
rect 737 2952 766 2957
rect 857 2957 862 2962
rect 857 2952 886 2957
rect 1521 2947 1526 2972
rect 1673 2962 1702 2967
rect 1729 2962 1782 2967
rect 1969 2962 2054 2967
rect 1969 2957 1974 2962
rect 177 2942 294 2947
rect 377 2942 470 2947
rect 601 2942 678 2947
rect 969 2942 1526 2947
rect 1537 2952 1558 2957
rect 1801 2952 1974 2957
rect 2049 2957 2054 2962
rect 2097 2957 2102 2972
rect 2049 2952 2102 2957
rect 2201 2957 2206 2972
rect 2249 2972 2382 2977
rect 2249 2957 2254 2972
rect 2201 2952 2254 2957
rect 2377 2957 2382 2972
rect 2377 2952 2406 2957
rect 969 2937 974 2942
rect 753 2932 974 2937
rect 753 2927 758 2932
rect 129 2922 222 2927
rect 217 2917 222 2922
rect 305 2922 366 2927
rect 505 2922 630 2927
rect 705 2922 758 2927
rect 1385 2922 1430 2927
rect 305 2917 310 2922
rect 217 2912 310 2917
rect 361 2907 366 2922
rect 705 2917 710 2922
rect 1425 2917 1430 2922
rect 1537 2917 1542 2952
rect 1721 2942 1774 2947
rect 1985 2942 2038 2947
rect 1985 2927 1990 2942
rect 2033 2937 2038 2942
rect 2113 2942 2198 2947
rect 2113 2937 2118 2942
rect 2033 2932 2118 2937
rect 2193 2937 2198 2942
rect 2281 2942 2334 2947
rect 2281 2937 2286 2942
rect 2193 2932 2286 2937
rect 2329 2937 2334 2942
rect 2417 2942 2790 2947
rect 2417 2937 2422 2942
rect 2329 2932 2422 2937
rect 1673 2922 1710 2927
rect 465 2912 710 2917
rect 729 2912 838 2917
rect 857 2912 1150 2917
rect 1345 2912 1374 2917
rect 1425 2912 1542 2917
rect 1705 2917 1710 2922
rect 1785 2922 1990 2927
rect 1785 2917 1790 2922
rect 1705 2912 1790 2917
rect 2017 2912 2054 2917
rect 2121 2912 2174 2917
rect 2441 2912 2502 2917
rect 465 2907 470 2912
rect 361 2902 470 2907
rect 617 2902 710 2907
rect 705 2897 710 2902
rect 817 2902 846 2907
rect 817 2897 822 2902
rect 705 2892 822 2897
rect 1329 2892 1406 2897
rect 1073 2882 1166 2887
rect 313 2872 438 2877
rect 897 2872 1046 2877
rect 1305 2872 1510 2877
rect 865 2852 934 2857
rect 1337 2842 1470 2847
rect 1489 2842 1630 2847
rect 1777 2842 1838 2847
rect 1449 2832 1478 2837
rect 2105 2832 2214 2837
rect 761 2822 918 2827
rect 1161 2822 1254 2827
rect 1369 2822 1430 2827
rect 1857 2822 1918 2827
rect 2233 2822 2342 2827
rect 2361 2822 2470 2827
rect 1641 2812 1686 2817
rect 1705 2812 1846 2817
rect 1841 2807 1846 2812
rect 1905 2812 2286 2817
rect 1905 2807 1910 2812
rect 945 2802 974 2807
rect 1209 2802 1310 2807
rect 1841 2802 1910 2807
rect 2281 2807 2286 2812
rect 2361 2812 2494 2817
rect 2361 2807 2366 2812
rect 2281 2802 2366 2807
rect 2745 2802 2822 2807
rect 2745 2797 2750 2802
rect 409 2792 470 2797
rect 529 2792 654 2797
rect 953 2792 1174 2797
rect 1441 2792 1486 2797
rect 1609 2792 1662 2797
rect 1753 2792 1790 2797
rect 1929 2792 2030 2797
rect 2721 2792 2750 2797
rect 2817 2797 2822 2802
rect 2817 2792 2846 2797
rect 529 2787 534 2792
rect 513 2782 534 2787
rect 649 2787 654 2792
rect 841 2787 934 2792
rect 1929 2787 1934 2792
rect 649 2782 678 2787
rect 817 2782 846 2787
rect 929 2782 974 2787
rect 1169 2782 1270 2787
rect 1585 2782 1614 2787
rect 513 2777 518 2782
rect 1609 2777 1614 2782
rect 1673 2782 1742 2787
rect 1673 2777 1678 2782
rect 433 2772 518 2777
rect 881 2772 1182 2777
rect 1353 2772 1582 2777
rect 1609 2772 1678 2777
rect 1737 2777 1742 2782
rect 1801 2782 1934 2787
rect 2025 2787 2030 2792
rect 2025 2782 2326 2787
rect 1801 2777 1806 2782
rect 2321 2777 2326 2782
rect 1737 2772 1806 2777
rect 1945 2772 2078 2777
rect 2321 2772 2854 2777
rect 433 2767 438 2772
rect 209 2762 438 2767
rect 577 2762 806 2767
rect 897 2762 1038 2767
rect 1465 2762 1550 2767
rect 2089 2762 2158 2767
rect 577 2757 582 2762
rect 897 2757 902 2762
rect 433 2752 582 2757
rect 593 2752 902 2757
rect 945 2752 1110 2757
rect 593 2747 598 2752
rect 201 2742 598 2747
rect 617 2742 790 2747
rect 1033 2742 1134 2747
rect 1145 2742 1254 2747
rect 1433 2742 1486 2747
rect 1761 2742 1806 2747
rect 2057 2742 2102 2747
rect 2217 2742 2286 2747
rect 2345 2742 2430 2747
rect 2633 2742 2694 2747
rect 2849 2742 2918 2747
rect 801 2737 918 2742
rect 1033 2737 1038 2742
rect 537 2732 574 2737
rect 593 2732 806 2737
rect 913 2732 1038 2737
rect 1057 2732 1118 2737
rect 1129 2732 1198 2737
rect 281 2727 422 2732
rect 593 2727 598 2732
rect 193 2722 286 2727
rect 417 2722 446 2727
rect 577 2722 598 2727
rect 665 2722 726 2727
rect 825 2722 894 2727
rect 281 2712 390 2717
rect 489 2712 550 2717
rect 641 2712 670 2717
rect 737 2712 878 2717
rect 961 2712 1046 2717
rect 665 2707 742 2712
rect 1057 2707 1062 2732
rect 1081 2722 1126 2727
rect 1393 2722 1558 2727
rect 2177 2722 2262 2727
rect 2761 2722 2894 2727
rect 2257 2717 2262 2722
rect 1113 2712 1198 2717
rect 1377 2712 1430 2717
rect 1641 2712 1686 2717
rect 1777 2712 1854 2717
rect 1873 2712 2046 2717
rect 2185 2712 2246 2717
rect 2257 2712 2374 2717
rect 2857 2712 2974 2717
rect 1777 2707 1782 2712
rect 529 2702 606 2707
rect 1057 2702 1166 2707
rect 1697 2702 1742 2707
rect 1753 2702 1782 2707
rect 1849 2707 1854 2712
rect 1849 2702 1886 2707
rect 2057 2702 2222 2707
rect 2713 2702 2758 2707
rect 737 2692 782 2697
rect 993 2692 1102 2697
rect 241 2682 310 2687
rect 377 2682 558 2687
rect 1729 2682 1790 2687
rect 1809 2682 1902 2687
rect 1937 2682 1990 2687
rect 2481 2682 2694 2687
rect 1633 2672 1710 2677
rect 2009 2672 2366 2677
rect 2385 2672 2446 2677
rect 1633 2667 1638 2672
rect 1705 2667 1790 2672
rect 1849 2667 2014 2672
rect 2361 2667 2366 2672
rect 913 2662 1078 2667
rect 1497 2662 1534 2667
rect 1609 2662 1638 2667
rect 1785 2662 1854 2667
rect 2361 2662 2414 2667
rect 913 2657 918 2662
rect 537 2652 582 2657
rect 889 2652 918 2657
rect 1073 2657 1078 2662
rect 2481 2657 2486 2682
rect 2689 2677 2694 2682
rect 2689 2672 2798 2677
rect 2793 2667 2798 2672
rect 2601 2662 2670 2667
rect 2793 2662 2822 2667
rect 2601 2657 2606 2662
rect 1073 2652 1102 2657
rect 1409 2652 1774 2657
rect 1865 2652 2486 2657
rect 2505 2652 2606 2657
rect 2665 2657 2670 2662
rect 2665 2652 2830 2657
rect 1769 2647 1870 2652
rect 1505 2642 1750 2647
rect 1889 2642 2566 2647
rect 2705 2642 2734 2647
rect 1889 2637 1894 2642
rect 2561 2637 2710 2642
rect 409 2632 470 2637
rect 553 2632 630 2637
rect 897 2632 934 2637
rect 993 2632 1094 2637
rect 1353 2632 1430 2637
rect 1449 2632 1894 2637
rect 1905 2632 2022 2637
rect 2129 2632 2350 2637
rect 2473 2632 2542 2637
rect 2345 2627 2478 2632
rect 377 2622 446 2627
rect 1441 2622 1630 2627
rect 1713 2622 1918 2627
rect 2097 2622 2326 2627
rect 2497 2622 2646 2627
rect 2657 2622 2878 2627
rect 1441 2617 1446 2622
rect 2657 2617 2662 2622
rect 585 2612 710 2617
rect 729 2612 782 2617
rect 1297 2612 1446 2617
rect 1457 2612 1486 2617
rect 2217 2612 2430 2617
rect 2625 2612 2662 2617
rect 585 2607 590 2612
rect 385 2602 590 2607
rect 705 2607 710 2612
rect 1457 2607 1462 2612
rect 1801 2607 1958 2612
rect 705 2602 878 2607
rect 1425 2602 1462 2607
rect 1745 2602 1806 2607
rect 1953 2602 2134 2607
rect 385 2597 390 2602
rect 2369 2597 2374 2612
rect 2505 2602 2742 2607
rect 153 2592 270 2597
rect 313 2592 390 2597
rect 545 2592 702 2597
rect 849 2592 950 2597
rect 1249 2592 1438 2597
rect 1465 2592 1566 2597
rect 1817 2592 1942 2597
rect 2369 2592 2398 2597
rect 2793 2592 2902 2597
rect 433 2582 518 2587
rect 769 2582 798 2587
rect 817 2582 1158 2587
rect 1417 2582 1630 2587
rect 1801 2582 1910 2587
rect 1961 2582 2038 2587
rect 2521 2582 2622 2587
rect 433 2577 438 2582
rect 305 2572 438 2577
rect 513 2577 518 2582
rect 1153 2577 1158 2582
rect 1961 2577 1966 2582
rect 513 2572 630 2577
rect 673 2572 878 2577
rect 969 2572 1078 2577
rect 1153 2572 1206 2577
rect 1353 2572 1382 2577
rect 1609 2572 1798 2577
rect 673 2567 678 2572
rect 873 2567 974 2572
rect 1377 2567 1534 2572
rect 1609 2567 1614 2572
rect 257 2562 678 2567
rect 697 2562 854 2567
rect 1529 2562 1614 2567
rect 1793 2567 1798 2572
rect 1897 2572 1966 2577
rect 2033 2577 2038 2582
rect 2033 2572 2542 2577
rect 1897 2567 1902 2572
rect 1793 2562 1902 2567
rect 1921 2562 2022 2567
rect 105 2552 398 2557
rect 393 2547 398 2552
rect 537 2552 726 2557
rect 537 2547 542 2552
rect 281 2542 334 2547
rect 393 2542 542 2547
rect 721 2547 726 2552
rect 801 2552 830 2557
rect 857 2552 974 2557
rect 1153 2552 1198 2557
rect 1361 2552 1510 2557
rect 1713 2552 1774 2557
rect 801 2547 806 2552
rect 721 2542 806 2547
rect 1097 2542 1150 2547
rect 1361 2537 1366 2552
rect 1505 2547 1510 2552
rect 1505 2542 1910 2547
rect 209 2532 286 2537
rect 945 2532 1086 2537
rect 1161 2532 1366 2537
rect 1905 2537 1910 2542
rect 2033 2542 2766 2547
rect 2033 2537 2038 2542
rect 1905 2532 2038 2537
rect 1081 2527 1166 2532
rect 1745 2522 1814 2527
rect 2953 2522 3080 2527
rect 1745 2517 1750 2522
rect 313 2512 374 2517
rect 393 2512 526 2517
rect 793 2512 934 2517
rect 1033 2512 1062 2517
rect 1057 2507 1062 2512
rect 1161 2512 1238 2517
rect 1441 2512 1478 2517
rect 1497 2512 1638 2517
rect 1721 2512 1750 2517
rect 1809 2517 1814 2522
rect 1809 2512 1838 2517
rect 2057 2512 2166 2517
rect 1161 2507 1166 2512
rect 1497 2507 1502 2512
rect 1057 2502 1166 2507
rect 1393 2502 1502 2507
rect 1633 2507 1638 2512
rect 1633 2502 1822 2507
rect 1889 2502 1958 2507
rect 1889 2497 1894 2502
rect 1185 2492 1326 2497
rect 1401 2492 1622 2497
rect 1617 2487 1622 2492
rect 1833 2492 1894 2497
rect 1953 2497 1958 2502
rect 1953 2492 2054 2497
rect 2689 2492 2830 2497
rect 1833 2487 1838 2492
rect 1385 2482 1558 2487
rect 1617 2482 1838 2487
rect 1009 2472 1214 2477
rect 1337 2472 1470 2477
rect 1497 2472 1526 2477
rect 1905 2472 1942 2477
rect 1937 2467 1942 2472
rect 2161 2472 2478 2477
rect 2161 2467 2166 2472
rect 1289 2462 1326 2467
rect 1321 2457 1326 2462
rect 1457 2462 1486 2467
rect 1577 2462 1886 2467
rect 1937 2462 1990 2467
rect 2137 2462 2166 2467
rect 2473 2467 2478 2472
rect 2473 2462 2502 2467
rect 1457 2457 1462 2462
rect 577 2452 662 2457
rect 577 2447 582 2452
rect 417 2442 582 2447
rect 657 2447 662 2452
rect 705 2452 990 2457
rect 1321 2452 1462 2457
rect 657 2442 686 2447
rect 705 2437 710 2452
rect 985 2447 990 2452
rect 1577 2447 1582 2462
rect 985 2442 1062 2447
rect 337 2432 446 2437
rect 649 2432 710 2437
rect 1057 2437 1062 2442
rect 1521 2442 1582 2447
rect 1881 2447 1886 2462
rect 2521 2452 2598 2457
rect 2521 2447 2526 2452
rect 1881 2442 1982 2447
rect 2009 2442 2118 2447
rect 2169 2442 2526 2447
rect 2593 2447 2598 2452
rect 2641 2452 2870 2457
rect 2641 2447 2646 2452
rect 2593 2442 2646 2447
rect 2865 2447 2870 2452
rect 2865 2442 2990 2447
rect 1521 2437 1526 2442
rect 2009 2437 2014 2442
rect 1057 2432 1526 2437
rect 1537 2432 1806 2437
rect 1865 2432 2014 2437
rect 2113 2437 2118 2442
rect 2113 2432 2142 2437
rect 2593 2432 2670 2437
rect 1537 2427 1542 2432
rect 2593 2427 2598 2432
rect 233 2422 286 2427
rect 593 2422 798 2427
rect 913 2422 998 2427
rect 1513 2422 1542 2427
rect 1601 2422 1646 2427
rect 1401 2417 1518 2422
rect 1953 2417 1958 2427
rect 2201 2422 2286 2427
rect 2329 2422 2414 2427
rect 2433 2422 2598 2427
rect 2609 2422 2782 2427
rect 2793 2422 2854 2427
rect 953 2412 1046 2417
rect 1041 2407 1046 2412
rect 1401 2407 1406 2417
rect 1809 2412 2318 2417
rect 1809 2407 1814 2412
rect 2313 2407 2318 2412
rect 2433 2407 2438 2422
rect 2897 2412 3080 2417
rect 417 2402 694 2407
rect 417 2397 422 2402
rect 97 2392 422 2397
rect 689 2397 694 2402
rect 737 2402 926 2407
rect 1041 2402 1102 2407
rect 1233 2402 1406 2407
rect 1425 2402 1582 2407
rect 1665 2402 1766 2407
rect 1785 2402 1814 2407
rect 1825 2402 1926 2407
rect 2193 2402 2294 2407
rect 2313 2402 2438 2407
rect 2473 2402 2542 2407
rect 2561 2402 2806 2407
rect 737 2397 742 2402
rect 689 2392 742 2397
rect 921 2397 926 2402
rect 1233 2397 1238 2402
rect 1665 2397 1670 2402
rect 921 2392 950 2397
rect 1121 2392 1238 2397
rect 1545 2392 1670 2397
rect 1761 2397 1766 2402
rect 2561 2397 2566 2402
rect 1761 2392 2182 2397
rect 2473 2392 2566 2397
rect 2801 2397 2806 2402
rect 2801 2392 2966 2397
rect 761 2387 894 2392
rect 1121 2387 1126 2392
rect 2177 2387 2182 2392
rect 249 2382 278 2387
rect 273 2367 278 2382
rect 433 2382 766 2387
rect 889 2382 1126 2387
rect 1953 2382 2038 2387
rect 2177 2382 2726 2387
rect 2921 2382 2950 2387
rect 433 2367 438 2382
rect 1761 2377 1854 2382
rect 2737 2377 2926 2382
rect 457 2372 486 2377
rect 713 2372 878 2377
rect 1593 2372 1766 2377
rect 1849 2372 1942 2377
rect 1985 2372 2030 2377
rect 2361 2372 2606 2377
rect 481 2367 718 2372
rect 1937 2367 1942 2372
rect 2209 2367 2342 2372
rect 2601 2367 2606 2372
rect 2689 2372 2742 2377
rect 2689 2367 2694 2372
rect 273 2362 438 2367
rect 865 2362 1302 2367
rect 1777 2362 1838 2367
rect 1937 2362 2214 2367
rect 2337 2362 2558 2367
rect 2601 2362 2694 2367
rect 2729 2362 2862 2367
rect 865 2357 870 2362
rect 513 2352 670 2357
rect 665 2347 670 2352
rect 809 2352 870 2357
rect 1377 2352 1446 2357
rect 1521 2352 1582 2357
rect 1729 2352 2006 2357
rect 2225 2352 2486 2357
rect 809 2347 814 2352
rect 1729 2347 1734 2352
rect 2481 2347 2486 2352
rect 2553 2352 2582 2357
rect 2881 2352 3054 2357
rect 2553 2347 2558 2352
rect 2881 2347 2886 2352
rect 497 2337 502 2347
rect 665 2342 814 2347
rect 1489 2342 1574 2347
rect 1633 2337 1638 2347
rect 1657 2342 1758 2347
rect 1769 2342 1790 2347
rect 2073 2342 2110 2347
rect 2241 2342 2358 2347
rect 2481 2342 2558 2347
rect 2673 2342 2886 2347
rect 3049 2347 3054 2352
rect 3049 2342 3080 2347
rect 497 2332 542 2337
rect 537 2327 542 2332
rect 617 2332 646 2337
rect 1361 2332 1390 2337
rect 1505 2332 1606 2337
rect 1633 2332 1686 2337
rect 617 2327 622 2332
rect 393 2322 518 2327
rect 537 2322 622 2327
rect 1385 2327 1390 2332
rect 1385 2322 1494 2327
rect 1489 2317 1494 2322
rect 1801 2322 2526 2327
rect 2785 2322 3080 2327
rect 1801 2317 1806 2322
rect 2785 2317 2790 2322
rect 1137 2312 1182 2317
rect 1489 2312 1806 2317
rect 1137 2307 1142 2312
rect 2001 2307 2006 2317
rect 2561 2312 2790 2317
rect 1057 2302 1142 2307
rect 1873 2302 1974 2307
rect 2001 2302 2478 2307
rect 2777 2302 2870 2307
rect 3049 2302 3080 2307
rect 3049 2297 3054 2302
rect 2457 2292 2550 2297
rect 2545 2287 2550 2292
rect 2897 2292 3054 2297
rect 377 2282 630 2287
rect 1569 2282 1926 2287
rect 2545 2282 2766 2287
rect 2761 2277 2766 2282
rect 2897 2277 2902 2292
rect 945 2272 1206 2277
rect 1433 2272 1550 2277
rect 2025 2272 2342 2277
rect 2761 2272 2902 2277
rect 1433 2267 1438 2272
rect 1257 2262 1326 2267
rect 1409 2262 1438 2267
rect 1545 2267 1550 2272
rect 1545 2262 1622 2267
rect 1257 2257 1262 2262
rect 65 2252 934 2257
rect 929 2247 934 2252
rect 1217 2252 1262 2257
rect 1321 2257 1326 2262
rect 1321 2252 1574 2257
rect 1217 2247 1222 2252
rect 929 2242 1222 2247
rect 1841 2242 1918 2247
rect 2353 2242 2406 2247
rect 1841 2237 1846 2242
rect 1273 2232 1310 2237
rect 1305 2227 1310 2232
rect 1457 2232 1558 2237
rect 1817 2232 1846 2237
rect 1913 2237 1918 2242
rect 1913 2232 1942 2237
rect 2617 2232 2702 2237
rect 1457 2227 1462 2232
rect 161 2222 326 2227
rect 793 2222 838 2227
rect 1305 2222 1462 2227
rect 1489 2222 1998 2227
rect 2217 2222 2382 2227
rect 2721 2222 2974 2227
rect 161 2217 166 2222
rect 0 2212 166 2217
rect 321 2217 326 2222
rect 2721 2217 2726 2222
rect 321 2212 350 2217
rect 921 2212 1014 2217
rect 1009 2207 1014 2212
rect 1033 2212 1254 2217
rect 1617 2212 1734 2217
rect 2201 2212 2238 2217
rect 2641 2212 2726 2217
rect 2969 2217 2974 2222
rect 2969 2212 3080 2217
rect 1033 2207 1038 2212
rect 1009 2202 1038 2207
rect 1249 2207 1254 2212
rect 1249 2202 1286 2207
rect 1713 2202 1822 2207
rect 2441 2202 2502 2207
rect 2649 2202 2678 2207
rect 0 2192 30 2197
rect 25 2187 30 2192
rect 177 2192 422 2197
rect 809 2192 886 2197
rect 905 2192 942 2197
rect 1009 2192 1014 2202
rect 2673 2197 2678 2202
rect 2737 2202 2790 2207
rect 2737 2197 2742 2202
rect 1721 2192 1750 2197
rect 177 2187 182 2192
rect 809 2187 814 2192
rect 25 2182 182 2187
rect 769 2182 814 2187
rect 881 2187 886 2192
rect 1241 2187 1310 2192
rect 1745 2187 1750 2192
rect 1825 2192 1854 2197
rect 1929 2192 2046 2197
rect 2081 2192 2438 2197
rect 2673 2192 2742 2197
rect 2825 2192 2958 2197
rect 1825 2187 1830 2192
rect 881 2182 1246 2187
rect 1305 2182 1398 2187
rect 1513 2182 1566 2187
rect 1745 2182 1830 2187
rect 2433 2177 2438 2192
rect 2521 2182 2630 2187
rect 2521 2177 2526 2182
rect 201 2172 270 2177
rect 1257 2172 1294 2177
rect 2433 2172 2526 2177
rect 2625 2177 2630 2182
rect 2625 2172 2886 2177
rect 2881 2167 2886 2172
rect 2953 2172 2982 2177
rect 2953 2167 2958 2172
rect 393 2162 478 2167
rect 825 2162 934 2167
rect 1609 2162 1846 2167
rect 2409 2162 2670 2167
rect 2881 2162 2958 2167
rect 1609 2157 1614 2162
rect 25 2152 182 2157
rect 25 2147 30 2152
rect 0 2142 30 2147
rect 177 2147 182 2152
rect 1025 2152 1134 2157
rect 1153 2152 1318 2157
rect 1553 2152 1614 2157
rect 1841 2157 1846 2162
rect 1841 2152 1870 2157
rect 2361 2152 2470 2157
rect 1025 2147 1030 2152
rect 177 2142 294 2147
rect 369 2142 470 2147
rect 793 2142 822 2147
rect 817 2137 822 2142
rect 897 2142 1030 2147
rect 1129 2147 1134 2152
rect 1129 2142 1302 2147
rect 1625 2142 1878 2147
rect 2113 2142 2166 2147
rect 2281 2142 2382 2147
rect 2489 2142 2606 2147
rect 2761 2142 2862 2147
rect 897 2137 902 2142
rect 2401 2137 2494 2142
rect 2601 2137 2606 2142
rect 817 2132 902 2137
rect 1257 2132 1310 2137
rect 1913 2132 1958 2137
rect 2289 2132 2406 2137
rect 2601 2132 2630 2137
rect 2737 2132 2782 2137
rect 1065 2127 1206 2132
rect 2801 2127 2918 2132
rect 0 2122 454 2127
rect 449 2117 454 2122
rect 489 2122 558 2127
rect 665 2122 782 2127
rect 1041 2122 1070 2127
rect 1201 2122 1230 2127
rect 489 2117 494 2122
rect 449 2112 494 2117
rect 553 2117 558 2122
rect 1225 2117 1230 2122
rect 1321 2122 1902 2127
rect 1321 2117 1326 2122
rect 553 2112 582 2117
rect 713 2112 742 2117
rect 937 2112 1022 2117
rect 1105 2112 1198 2117
rect 1225 2112 1326 2117
rect 1897 2117 1902 2122
rect 1969 2122 2054 2127
rect 2201 2122 2806 2127
rect 2913 2122 3080 2127
rect 1969 2117 1974 2122
rect 1897 2112 1974 2117
rect 2113 2112 2222 2117
rect 2329 2112 2438 2117
rect 2729 2112 2774 2117
rect 2817 2112 2902 2117
rect 937 2107 942 2112
rect 0 2102 30 2107
rect 25 2097 30 2102
rect 217 2102 446 2107
rect 601 2102 678 2107
rect 729 2102 942 2107
rect 1017 2107 1022 2112
rect 1665 2107 1782 2112
rect 1017 2102 1046 2107
rect 217 2097 222 2102
rect 601 2097 606 2102
rect 25 2092 222 2097
rect 433 2092 486 2097
rect 537 2092 606 2097
rect 673 2097 678 2102
rect 1041 2097 1046 2102
rect 1105 2102 1134 2107
rect 1513 2102 1670 2107
rect 1777 2102 1806 2107
rect 2425 2102 2518 2107
rect 2585 2102 2814 2107
rect 1105 2097 1110 2102
rect 2809 2097 2814 2102
rect 3049 2102 3080 2107
rect 3049 2097 3054 2102
rect 673 2092 822 2097
rect 953 2092 990 2097
rect 1041 2092 1110 2097
rect 1169 2092 1206 2097
rect 1649 2092 1750 2097
rect 1825 2092 2054 2097
rect 2721 2092 2790 2097
rect 2809 2092 3054 2097
rect 1825 2087 1830 2092
rect 449 2082 766 2087
rect 969 2082 1022 2087
rect 1697 2082 1830 2087
rect 2049 2087 2054 2092
rect 2049 2082 2174 2087
rect 2353 2082 2758 2087
rect 241 2072 374 2077
rect 393 2072 734 2077
rect 2137 2072 2198 2077
rect 2273 2072 2390 2077
rect 241 2067 246 2072
rect 0 2062 246 2067
rect 369 2067 374 2072
rect 2385 2067 2390 2072
rect 2753 2072 2782 2077
rect 2753 2067 2758 2072
rect 369 2062 398 2067
rect 497 2062 678 2067
rect 1097 2062 1262 2067
rect 1737 2062 2038 2067
rect 2289 2062 2366 2067
rect 2385 2062 2758 2067
rect 393 2057 502 2062
rect 521 2047 630 2052
rect 1097 2047 1102 2062
rect 257 2042 526 2047
rect 625 2042 654 2047
rect 1017 2042 1102 2047
rect 1257 2047 1262 2062
rect 1257 2042 1286 2047
rect 1833 2042 2166 2047
rect 2873 2042 2998 2047
rect 401 2032 430 2037
rect 537 2032 646 2037
rect 1113 2032 1198 2037
rect 1225 2032 1318 2037
rect 1369 2032 1438 2037
rect 1625 2032 1734 2037
rect 2337 2032 2446 2037
rect 2617 2032 2742 2037
rect 2761 2032 2870 2037
rect 425 2027 542 2032
rect 641 2017 646 2032
rect 1313 2027 1318 2032
rect 1073 2022 1166 2027
rect 1257 2022 1302 2027
rect 1313 2022 1406 2027
rect 1753 2022 1966 2027
rect 2185 2022 2238 2027
rect 1625 2017 1758 2022
rect 1961 2017 1966 2022
rect 2617 2017 2622 2032
rect 0 2012 238 2017
rect 313 2012 422 2017
rect 513 2012 606 2017
rect 641 2012 726 2017
rect 953 2012 1006 2017
rect 1601 2012 1630 2017
rect 1961 2012 1990 2017
rect 2009 2012 2166 2017
rect 2593 2012 2622 2017
rect 2737 2017 2742 2032
rect 2737 2012 3080 2017
rect 1777 2007 1942 2012
rect 2009 2007 2014 2012
rect 2161 2007 2246 2012
rect 809 2002 918 2007
rect 1281 2002 1478 2007
rect 1489 2002 1782 2007
rect 1937 2002 2014 2007
rect 2241 2002 2766 2007
rect 505 1992 534 1997
rect 529 1987 534 1992
rect 633 1992 886 1997
rect 937 1992 1182 1997
rect 1569 1992 1630 1997
rect 1705 1992 1894 1997
rect 1905 1992 1966 1997
rect 2025 1992 2230 1997
rect 633 1987 638 1992
rect 529 1982 638 1987
rect 881 1987 886 1992
rect 2225 1987 2230 1992
rect 2409 1992 2438 1997
rect 2625 1992 2806 1997
rect 2865 1992 2942 1997
rect 2409 1987 2414 1992
rect 881 1982 910 1987
rect 905 1977 910 1982
rect 993 1982 1102 1987
rect 1665 1982 1694 1987
rect 1785 1982 1846 1987
rect 2225 1982 2414 1987
rect 2673 1982 2726 1987
rect 993 1977 998 1982
rect 1121 1977 1190 1982
rect 1689 1977 1790 1982
rect 905 1972 998 1977
rect 1073 1972 1126 1977
rect 1185 1972 1382 1977
rect 2625 1972 2918 1977
rect 657 1962 886 1967
rect 1017 1962 1174 1967
rect 1657 1962 1742 1967
rect 1657 1957 1662 1962
rect 353 1952 446 1957
rect 1033 1952 1062 1957
rect 353 1947 358 1952
rect 201 1942 230 1947
rect 329 1942 358 1947
rect 441 1947 446 1952
rect 1057 1947 1062 1952
rect 1121 1952 1318 1957
rect 1561 1952 1662 1957
rect 1737 1957 1742 1962
rect 1801 1962 2014 1967
rect 1801 1957 1806 1962
rect 1737 1952 1806 1957
rect 2009 1957 2014 1962
rect 2073 1962 2238 1967
rect 2305 1962 2590 1967
rect 2705 1962 2774 1967
rect 2073 1957 2078 1962
rect 2009 1952 2078 1957
rect 2233 1957 2238 1962
rect 2233 1952 2262 1957
rect 2673 1952 2758 1957
rect 2881 1952 2982 1957
rect 1121 1947 1126 1952
rect 441 1942 470 1947
rect 825 1942 958 1947
rect 1057 1942 1126 1947
rect 1145 1942 1182 1947
rect 1257 1942 1310 1947
rect 1617 1942 1726 1947
rect 1817 1942 1982 1947
rect 2089 1942 2230 1947
rect 2353 1942 2374 1947
rect 2417 1942 2462 1947
rect 2729 1942 2766 1947
rect 2225 1937 2310 1942
rect 1225 1932 1398 1937
rect 1577 1932 1806 1937
rect 1969 1932 1998 1937
rect 1801 1927 1974 1932
rect 2305 1927 2310 1937
rect 321 1922 510 1927
rect 617 1922 934 1927
rect 961 1922 1062 1927
rect 1217 1922 1254 1927
rect 1297 1922 1326 1927
rect 2305 1922 2358 1927
rect 433 1912 510 1917
rect 833 1912 838 1922
rect 2369 1917 2374 1942
rect 2953 1922 3080 1927
rect 1081 1912 1246 1917
rect 1769 1912 2374 1917
rect 2409 1912 2566 1917
rect 1217 1902 1414 1907
rect 1113 1897 1190 1902
rect 297 1892 1118 1897
rect 1185 1892 1214 1897
rect 1129 1882 1190 1887
rect 1209 1877 1214 1892
rect 1425 1892 1486 1897
rect 2249 1892 2278 1897
rect 1425 1877 1430 1892
rect 2273 1887 2278 1892
rect 2369 1892 2398 1897
rect 2369 1887 2374 1892
rect 1849 1882 1902 1887
rect 2017 1882 2166 1887
rect 2273 1882 2374 1887
rect 249 1872 382 1877
rect 497 1872 590 1877
rect 793 1872 1134 1877
rect 1209 1872 1430 1877
rect 2425 1872 2646 1877
rect 249 1862 278 1867
rect 393 1862 510 1867
rect 601 1862 766 1867
rect 273 1857 398 1862
rect 505 1857 606 1862
rect 2425 1857 2430 1872
rect 913 1852 1030 1857
rect 2097 1852 2126 1857
rect 2345 1852 2430 1857
rect 2641 1857 2646 1872
rect 2641 1852 2774 1857
rect 913 1847 918 1852
rect 129 1842 918 1847
rect 1025 1847 1030 1852
rect 1025 1842 1510 1847
rect 1977 1842 2078 1847
rect 2097 1842 2158 1847
rect 2441 1842 2630 1847
rect 2977 1842 3054 1847
rect 1977 1837 1982 1842
rect 929 1832 1014 1837
rect 1865 1832 1934 1837
rect 1953 1832 1982 1837
rect 2073 1837 2078 1842
rect 2073 1832 2190 1837
rect 2209 1832 2310 1837
rect 2329 1832 2438 1837
rect 929 1827 934 1832
rect 2209 1827 2214 1832
rect 281 1822 326 1827
rect 449 1822 934 1827
rect 945 1817 950 1827
rect 1201 1822 1334 1827
rect 1369 1822 1422 1827
rect 1697 1822 1846 1827
rect 1953 1822 2214 1827
rect 2305 1827 2310 1832
rect 2305 1822 2726 1827
rect 2769 1822 2822 1827
rect 2857 1822 2902 1827
rect 0 1812 174 1817
rect 537 1812 566 1817
rect 945 1812 1190 1817
rect 1249 1812 1278 1817
rect 401 1807 470 1812
rect 1185 1807 1254 1812
rect 1697 1807 1702 1822
rect 1841 1817 1846 1822
rect 2977 1817 2982 1842
rect 3049 1837 3054 1842
rect 3049 1832 3080 1837
rect 1841 1812 1934 1817
rect 2241 1812 2430 1817
rect 2913 1812 2982 1817
rect 3009 1817 3014 1827
rect 3009 1812 3080 1817
rect 201 1802 406 1807
rect 465 1802 494 1807
rect 641 1802 750 1807
rect 1273 1802 1310 1807
rect 1545 1802 1638 1807
rect 1673 1802 1702 1807
rect 1929 1807 1934 1812
rect 2073 1807 2206 1812
rect 2601 1807 2742 1812
rect 2913 1807 2918 1812
rect 1929 1802 2078 1807
rect 2201 1802 2230 1807
rect 2577 1802 2606 1807
rect 2737 1802 2918 1807
rect 513 1797 622 1802
rect 2225 1797 2230 1802
rect 2249 1797 2510 1802
rect 97 1792 134 1797
rect 417 1792 518 1797
rect 617 1792 894 1797
rect 1145 1792 1254 1797
rect 1145 1787 1150 1792
rect 369 1782 558 1787
rect 617 1782 678 1787
rect 857 1782 1038 1787
rect 1097 1782 1150 1787
rect 1249 1787 1254 1792
rect 1329 1792 1414 1797
rect 1465 1792 1550 1797
rect 1329 1787 1334 1792
rect 1249 1782 1334 1787
rect 1409 1787 1414 1792
rect 1545 1787 1550 1792
rect 1657 1792 1918 1797
rect 2089 1792 2214 1797
rect 2225 1792 2254 1797
rect 2505 1792 2670 1797
rect 2705 1792 2726 1797
rect 3049 1792 3080 1797
rect 1657 1787 1662 1792
rect 1913 1787 2094 1792
rect 2209 1787 2214 1792
rect 3049 1787 3054 1792
rect 1409 1782 1430 1787
rect 1425 1777 1430 1782
rect 1497 1782 1526 1787
rect 1545 1782 1662 1787
rect 2209 1782 2494 1787
rect 2641 1782 2734 1787
rect 2753 1782 2854 1787
rect 1497 1777 1502 1782
rect 2753 1777 2758 1782
rect 0 1772 86 1777
rect 81 1767 86 1772
rect 145 1772 358 1777
rect 545 1772 598 1777
rect 145 1767 150 1772
rect 353 1767 454 1772
rect 545 1767 550 1772
rect 81 1762 150 1767
rect 449 1762 550 1767
rect 593 1767 598 1772
rect 657 1772 686 1777
rect 1161 1772 1286 1777
rect 1425 1772 1502 1777
rect 1721 1772 2758 1777
rect 2849 1777 2854 1782
rect 2913 1782 3054 1787
rect 2849 1772 2878 1777
rect 657 1767 662 1772
rect 2913 1767 2918 1782
rect 593 1762 662 1767
rect 713 1762 1214 1767
rect 1297 1762 1398 1767
rect 1681 1762 1710 1767
rect 2065 1762 2326 1767
rect 2345 1762 2478 1767
rect 2673 1762 2918 1767
rect 1209 1757 1302 1762
rect 1705 1757 2070 1762
rect 2673 1757 2678 1762
rect 369 1752 422 1757
rect 1097 1752 1190 1757
rect 2089 1752 2182 1757
rect 2465 1752 2678 1757
rect 2697 1752 2766 1757
rect 369 1747 374 1752
rect 1185 1747 1190 1752
rect 2177 1747 2182 1752
rect 2281 1747 2470 1752
rect 321 1742 374 1747
rect 393 1742 430 1747
rect 753 1742 854 1747
rect 865 1742 966 1747
rect 1033 1742 1110 1747
rect 1185 1742 1390 1747
rect 1521 1742 1726 1747
rect 849 1737 854 1742
rect 1721 1737 1726 1742
rect 1785 1742 2030 1747
rect 2177 1742 2286 1747
rect 2489 1742 2534 1747
rect 2657 1742 2750 1747
rect 2857 1742 2902 1747
rect 2977 1742 3062 1747
rect 1785 1737 1790 1742
rect 2977 1737 2982 1742
rect 545 1732 798 1737
rect 849 1732 878 1737
rect 1001 1732 1030 1737
rect 1113 1732 1182 1737
rect 1721 1732 1790 1737
rect 2073 1732 2158 1737
rect 2305 1732 2430 1737
rect 2953 1732 2982 1737
rect 3057 1737 3062 1742
rect 3057 1732 3080 1737
rect 545 1727 550 1732
rect 873 1727 1006 1732
rect 0 1722 310 1727
rect 305 1717 310 1722
rect 377 1722 550 1727
rect 785 1722 854 1727
rect 1249 1722 1286 1727
rect 1649 1722 1702 1727
rect 1921 1722 2038 1727
rect 377 1717 382 1722
rect 849 1717 854 1722
rect 1921 1717 1926 1722
rect 305 1712 382 1717
rect 761 1712 806 1717
rect 849 1712 1054 1717
rect 1897 1712 1926 1717
rect 2033 1717 2038 1722
rect 2177 1722 2286 1727
rect 2609 1722 2694 1727
rect 3075 1722 3080 1732
rect 2177 1717 2182 1722
rect 2033 1712 2182 1717
rect 2281 1717 2286 1722
rect 2281 1712 3078 1717
rect 1785 1702 1894 1707
rect 1945 1702 2022 1707
rect 2233 1702 2270 1707
rect 2569 1702 2598 1707
rect 2697 1702 2790 1707
rect 2593 1697 2702 1702
rect 401 1692 494 1697
rect 905 1692 1142 1697
rect 1945 1692 2222 1697
rect 2281 1692 2462 1697
rect 2217 1687 2286 1692
rect 3075 1687 3080 1707
rect 817 1682 886 1687
rect 1953 1682 2046 1687
rect 2497 1682 2574 1687
rect 2593 1682 3080 1687
rect 817 1677 822 1682
rect 881 1677 966 1682
rect 2497 1677 2502 1682
rect 425 1672 566 1677
rect 793 1672 822 1677
rect 961 1672 1222 1677
rect 1265 1672 1414 1677
rect 2185 1672 2502 1677
rect 2569 1677 2574 1682
rect 2569 1672 2662 1677
rect 897 1662 950 1667
rect 1265 1657 1270 1672
rect 617 1652 662 1657
rect 809 1652 886 1657
rect 1001 1652 1166 1657
rect 1209 1652 1270 1657
rect 1409 1657 1414 1672
rect 1665 1662 1942 1667
rect 1937 1657 1942 1662
rect 2025 1662 2126 1667
rect 2513 1662 2718 1667
rect 2025 1657 2030 1662
rect 2313 1657 2398 1662
rect 1409 1652 1678 1657
rect 1937 1652 2030 1657
rect 2289 1652 2318 1657
rect 2393 1652 2486 1657
rect 1001 1647 1006 1652
rect 273 1642 398 1647
rect 473 1642 606 1647
rect 673 1642 750 1647
rect 865 1642 1006 1647
rect 1161 1647 1166 1652
rect 2513 1647 2518 1662
rect 2537 1652 2774 1657
rect 2769 1647 2774 1652
rect 1161 1642 1190 1647
rect 1281 1642 1398 1647
rect 2137 1642 2382 1647
rect 2489 1642 2518 1647
rect 2641 1642 2670 1647
rect 2769 1642 2966 1647
rect 2985 1642 3054 1647
rect 273 1627 278 1642
rect 393 1637 398 1642
rect 601 1637 678 1642
rect 2377 1637 2494 1642
rect 2665 1637 2758 1642
rect 2985 1637 2990 1642
rect 393 1632 422 1637
rect 993 1632 1150 1637
rect 2753 1632 2782 1637
rect 2961 1632 2990 1637
rect 3049 1637 3054 1642
rect 3049 1632 3080 1637
rect 193 1622 278 1627
rect 345 1622 454 1627
rect 489 1622 1126 1627
rect 1201 1622 1462 1627
rect 1681 1622 1758 1627
rect 1921 1622 1998 1627
rect 2201 1622 2246 1627
rect 2265 1622 2758 1627
rect 1921 1617 1926 1622
rect 2753 1617 2758 1622
rect 257 1612 286 1617
rect 857 1612 1262 1617
rect 1545 1612 1614 1617
rect 1737 1612 1926 1617
rect 1961 1612 2006 1617
rect 2113 1612 2182 1617
rect 2513 1612 2542 1617
rect 2753 1612 3080 1617
rect 2113 1607 2118 1612
rect 649 1602 774 1607
rect 929 1602 1102 1607
rect 1273 1602 1382 1607
rect 1545 1602 1606 1607
rect 2089 1602 2118 1607
rect 2177 1607 2182 1612
rect 2441 1607 2518 1612
rect 2177 1602 2254 1607
rect 2297 1602 2446 1607
rect 2633 1602 2758 1607
rect 1097 1597 1278 1602
rect 2753 1597 2758 1602
rect 585 1592 750 1597
rect 825 1592 886 1597
rect 1001 1592 1078 1597
rect 1633 1592 1862 1597
rect 2017 1592 2158 1597
rect 2457 1592 2486 1597
rect 2753 1592 2846 1597
rect 633 1582 742 1587
rect 809 1582 894 1587
rect 1113 1582 1286 1587
rect 1281 1577 1286 1582
rect 1361 1582 1390 1587
rect 1633 1582 1638 1592
rect 2153 1587 2462 1592
rect 2841 1587 2846 1592
rect 2953 1592 3080 1597
rect 2953 1587 2958 1592
rect 1985 1582 2134 1587
rect 2513 1582 2686 1587
rect 2841 1582 2958 1587
rect 1361 1577 1366 1582
rect 2513 1577 2518 1582
rect 753 1567 758 1577
rect 1033 1572 1126 1577
rect 1281 1572 1366 1577
rect 1465 1572 1974 1577
rect 2145 1572 2222 1577
rect 2273 1572 2470 1577
rect 2489 1572 2518 1577
rect 2681 1577 2686 1582
rect 2681 1572 2822 1577
rect 1969 1567 2150 1572
rect 2273 1567 2278 1572
rect 753 1562 1150 1567
rect 1649 1562 1702 1567
rect 2249 1562 2278 1567
rect 2465 1567 2470 1572
rect 2465 1562 2670 1567
rect 2977 1562 3080 1567
rect 569 1552 734 1557
rect 1025 1552 1158 1557
rect 1177 1552 1262 1557
rect 1713 1552 1846 1557
rect 2017 1552 2110 1557
rect 2257 1552 2494 1557
rect 2841 1552 2958 1557
rect 569 1547 574 1552
rect 257 1542 574 1547
rect 729 1547 734 1552
rect 817 1547 886 1552
rect 1177 1547 1182 1552
rect 729 1542 822 1547
rect 881 1542 910 1547
rect 1097 1542 1182 1547
rect 1257 1547 1262 1552
rect 2841 1547 2846 1552
rect 1257 1542 1318 1547
rect 1737 1542 1766 1547
rect 1761 1537 1766 1542
rect 1825 1542 1998 1547
rect 2129 1542 2230 1547
rect 1825 1537 1830 1542
rect 1993 1537 2134 1542
rect 2225 1537 2230 1542
rect 2257 1542 2294 1547
rect 2401 1542 2846 1547
rect 2953 1547 2958 1552
rect 2953 1542 3080 1547
rect 2257 1537 2262 1542
rect 513 1532 742 1537
rect 833 1532 862 1537
rect 1761 1532 1830 1537
rect 2225 1532 2262 1537
rect 0 1522 150 1527
rect 241 1522 326 1527
rect 145 1517 150 1522
rect 321 1517 326 1522
rect 513 1517 518 1532
rect 737 1527 838 1532
rect 1057 1527 1190 1532
rect 2281 1527 2854 1532
rect 2977 1527 2982 1537
rect 529 1522 606 1527
rect 689 1522 718 1527
rect 145 1512 222 1517
rect 321 1512 518 1517
rect 713 1517 718 1522
rect 873 1522 1062 1527
rect 1185 1522 1246 1527
rect 1905 1522 2286 1527
rect 2849 1522 2982 1527
rect 2993 1522 3080 1527
rect 873 1517 878 1522
rect 1905 1517 1910 1522
rect 2993 1517 2998 1522
rect 713 1512 878 1517
rect 1073 1512 1174 1517
rect 1505 1512 1678 1517
rect 1849 1512 1910 1517
rect 1953 1512 2838 1517
rect 2833 1507 2838 1512
rect 2969 1512 2998 1517
rect 2969 1507 2974 1512
rect 233 1502 286 1507
rect 601 1502 678 1507
rect 673 1497 678 1502
rect 905 1502 950 1507
rect 1209 1502 1254 1507
rect 1345 1502 1390 1507
rect 2089 1502 2326 1507
rect 2473 1502 2654 1507
rect 2777 1502 2814 1507
rect 2833 1502 2974 1507
rect 2993 1502 3080 1507
rect 905 1497 910 1502
rect 2321 1497 2478 1502
rect 673 1492 910 1497
rect 2057 1492 2134 1497
rect 2225 1492 2254 1497
rect 2273 1492 2302 1497
rect 2129 1487 2230 1492
rect 2297 1487 2302 1492
rect 2521 1492 2598 1497
rect 2521 1487 2526 1492
rect 2297 1482 2526 1487
rect 2593 1487 2598 1492
rect 2593 1482 2790 1487
rect 2785 1477 2790 1482
rect 2833 1482 2982 1487
rect 2833 1477 2838 1482
rect 289 1472 494 1477
rect 577 1472 638 1477
rect 1049 1472 1254 1477
rect 2105 1472 2206 1477
rect 857 1462 1006 1467
rect 0 1452 174 1457
rect 729 1452 822 1457
rect 729 1447 734 1452
rect 257 1442 734 1447
rect 817 1437 822 1452
rect 857 1447 862 1462
rect 833 1442 862 1447
rect 1001 1447 1006 1462
rect 1049 1457 1054 1472
rect 1025 1452 1054 1457
rect 1249 1457 1254 1472
rect 2201 1467 2206 1472
rect 2545 1472 2574 1477
rect 2785 1472 2838 1477
rect 2977 1477 2982 1482
rect 2993 1477 2998 1502
rect 3009 1482 3080 1487
rect 2977 1472 2998 1477
rect 2545 1467 2550 1472
rect 1297 1462 1382 1467
rect 1865 1462 2182 1467
rect 2201 1462 2550 1467
rect 2737 1457 2878 1462
rect 1249 1452 1358 1457
rect 2657 1452 2742 1457
rect 2873 1452 2966 1457
rect 1001 1442 1230 1447
rect 1265 1442 1310 1447
rect 2753 1442 2862 1447
rect 129 1432 230 1437
rect 657 1432 798 1437
rect 817 1432 998 1437
rect 1185 1432 1222 1437
rect 1585 1432 1654 1437
rect 1713 1432 1742 1437
rect 1585 1427 1590 1432
rect 321 1422 622 1427
rect 753 1422 838 1427
rect 945 1422 1006 1427
rect 1081 1422 1126 1427
rect 1233 1422 1390 1427
rect 1561 1422 1590 1427
rect 1649 1427 1654 1432
rect 1649 1422 1678 1427
rect 1705 1422 1766 1427
rect 2017 1422 2118 1427
rect 2321 1422 2918 1427
rect 321 1402 326 1422
rect 2913 1417 2918 1422
rect 737 1412 782 1417
rect 1585 1412 1750 1417
rect 1937 1412 1974 1417
rect 2913 1412 3080 1417
rect 1265 1407 1334 1412
rect 433 1402 742 1407
rect 1009 1402 1094 1407
rect 1137 1402 1270 1407
rect 1329 1402 1430 1407
rect 1457 1402 1846 1407
rect 185 1392 342 1397
rect 745 1392 854 1397
rect 865 1392 1038 1397
rect 1281 1392 1318 1397
rect 1561 1392 1614 1397
rect 1673 1392 1958 1397
rect 1993 1392 2190 1397
rect 2289 1392 2478 1397
rect 2609 1392 2934 1397
rect 865 1387 870 1392
rect 1313 1387 1318 1392
rect 1993 1387 1998 1392
rect 617 1382 870 1387
rect 1169 1382 1302 1387
rect 1313 1382 1446 1387
rect 1617 1382 1862 1387
rect 1873 1382 1998 1387
rect 2185 1387 2190 1392
rect 2185 1382 2262 1387
rect 1857 1377 1862 1382
rect 2257 1377 2374 1382
rect 449 1372 518 1377
rect 625 1372 654 1377
rect 865 1372 982 1377
rect 1529 1372 1790 1377
rect 1857 1372 2054 1377
rect 2369 1372 2614 1377
rect 649 1367 870 1372
rect 1441 1367 1510 1372
rect 2169 1367 2238 1372
rect 1153 1362 1222 1367
rect 1369 1362 1446 1367
rect 1505 1362 2006 1367
rect 2065 1362 2174 1367
rect 2233 1362 2558 1367
rect 2745 1362 2902 1367
rect 2921 1362 2982 1367
rect 2001 1357 2070 1362
rect 137 1352 1142 1357
rect 1137 1347 1142 1352
rect 1225 1352 1358 1357
rect 1457 1352 1550 1357
rect 1225 1347 1230 1352
rect 1353 1347 1462 1352
rect 1545 1347 1550 1352
rect 1641 1352 1670 1357
rect 1769 1352 1814 1357
rect 1897 1352 1982 1357
rect 2185 1352 2222 1357
rect 2321 1352 2350 1357
rect 2457 1352 2502 1357
rect 1641 1347 1646 1352
rect 1809 1347 1902 1352
rect 2217 1347 2310 1352
rect 1137 1342 1230 1347
rect 1481 1342 1526 1347
rect 1545 1342 1646 1347
rect 1697 1342 1790 1347
rect 417 1332 470 1337
rect 729 1332 814 1337
rect 825 1332 950 1337
rect 1249 1332 1342 1337
rect 1249 1327 1254 1332
rect 0 1322 302 1327
rect 433 1322 790 1327
rect 897 1322 990 1327
rect 1121 1322 1254 1327
rect 1337 1327 1342 1332
rect 1385 1332 1454 1337
rect 1385 1327 1390 1332
rect 1337 1322 1390 1327
rect 1449 1327 1454 1332
rect 1521 1327 1526 1342
rect 1697 1327 1702 1342
rect 1785 1337 1790 1342
rect 1921 1342 2198 1347
rect 2305 1342 2398 1347
rect 1921 1337 1926 1342
rect 2393 1337 2398 1342
rect 2489 1342 2518 1347
rect 2545 1342 2726 1347
rect 2489 1337 2494 1342
rect 1761 1327 1766 1337
rect 1785 1332 1926 1337
rect 1945 1332 2022 1337
rect 2257 1332 2334 1337
rect 2393 1332 2494 1337
rect 1449 1322 1478 1327
rect 1521 1322 1702 1327
rect 1721 1322 1766 1327
rect 1985 1322 2038 1327
rect 2561 1322 2670 1327
rect 2761 1322 2806 1327
rect 2561 1317 2566 1322
rect 265 1312 350 1317
rect 673 1312 790 1317
rect 785 1307 790 1312
rect 881 1312 910 1317
rect 1065 1312 1182 1317
rect 1265 1312 1374 1317
rect 1433 1312 1502 1317
rect 2017 1312 2126 1317
rect 2161 1312 2374 1317
rect 2537 1312 2566 1317
rect 2665 1317 2670 1322
rect 2801 1317 2806 1322
rect 2665 1312 2766 1317
rect 2801 1312 2822 1317
rect 881 1307 886 1312
rect 425 1302 462 1307
rect 785 1302 886 1307
rect 1001 1302 1086 1307
rect 1777 1302 1862 1307
rect 2049 1302 2094 1307
rect 265 1292 294 1297
rect 2089 1287 2094 1302
rect 2353 1302 2446 1307
rect 2561 1302 2654 1307
rect 2353 1297 2358 1302
rect 2273 1292 2358 1297
rect 2753 1292 2878 1297
rect 2273 1287 2278 1292
rect 929 1282 990 1287
rect 985 1277 990 1282
rect 1097 1282 1422 1287
rect 2089 1282 2278 1287
rect 2377 1282 2486 1287
rect 1097 1277 1102 1282
rect 2377 1277 2382 1282
rect 985 1272 1102 1277
rect 1441 1272 1518 1277
rect 2297 1272 2382 1277
rect 2481 1277 2486 1282
rect 2481 1272 2726 1277
rect 2745 1272 2846 1277
rect 1377 1267 1446 1272
rect 1513 1267 1518 1272
rect 2721 1267 2726 1272
rect 1313 1262 1382 1267
rect 1513 1262 1974 1267
rect 2337 1262 2486 1267
rect 2721 1262 2998 1267
rect 2521 1257 2702 1262
rect 353 1252 790 1257
rect 1233 1252 1302 1257
rect 353 1247 358 1252
rect 249 1242 358 1247
rect 785 1247 790 1252
rect 1297 1247 1302 1252
rect 1457 1252 1502 1257
rect 2441 1252 2526 1257
rect 2697 1252 2782 1257
rect 1457 1247 1462 1252
rect 785 1242 1086 1247
rect 1297 1242 1462 1247
rect 2097 1242 2310 1247
rect 2361 1242 2430 1247
rect 2497 1242 2526 1247
rect 2545 1242 2702 1247
rect 2753 1242 2854 1247
rect 2097 1237 2102 1242
rect 2425 1237 2502 1242
rect 1697 1232 1822 1237
rect 1857 1232 2102 1237
rect 2297 1232 2350 1237
rect 2553 1232 2582 1237
rect 2737 1232 2766 1237
rect 2857 1232 2942 1237
rect 2577 1227 2742 1232
rect 153 1222 302 1227
rect 369 1222 454 1227
rect 465 1222 710 1227
rect 737 1222 774 1227
rect 985 1222 1134 1227
rect 1417 1222 1654 1227
rect 2441 1222 2542 1227
rect 737 1217 742 1222
rect 241 1212 294 1217
rect 689 1212 742 1217
rect 793 1212 942 1217
rect 1273 1212 1406 1217
rect 2193 1212 2430 1217
rect 2553 1212 3080 1217
rect 313 1202 422 1207
rect 441 1202 550 1207
rect 569 1202 670 1207
rect 313 1197 318 1202
rect 169 1192 318 1197
rect 417 1197 422 1202
rect 569 1197 574 1202
rect 665 1197 742 1202
rect 793 1197 798 1212
rect 417 1192 574 1197
rect 737 1192 798 1197
rect 937 1197 942 1212
rect 2425 1207 2558 1212
rect 1041 1202 1214 1207
rect 1481 1202 1630 1207
rect 937 1192 966 1197
rect 1185 1192 1294 1197
rect 1377 1192 1462 1197
rect 1481 1187 1486 1202
rect 105 1182 158 1187
rect 153 1167 158 1182
rect 297 1182 438 1187
rect 489 1182 726 1187
rect 809 1182 1006 1187
rect 1233 1182 1486 1187
rect 1625 1187 1630 1202
rect 1793 1202 2126 1207
rect 1689 1192 1774 1197
rect 1793 1187 1798 1202
rect 2121 1187 2126 1202
rect 2289 1192 2414 1197
rect 2425 1192 2550 1197
rect 2873 1192 2902 1197
rect 2897 1187 2902 1192
rect 2969 1192 2998 1197
rect 2969 1187 2974 1192
rect 1625 1182 1646 1187
rect 297 1167 302 1182
rect 721 1177 814 1182
rect 1641 1177 1646 1182
rect 1721 1182 1798 1187
rect 2009 1182 2086 1187
rect 2121 1182 2534 1187
rect 2569 1182 2734 1187
rect 2897 1182 2974 1187
rect 1721 1177 1726 1182
rect 2009 1177 2014 1182
rect 529 1172 702 1177
rect 1001 1172 1286 1177
rect 1281 1167 1286 1172
rect 1417 1172 1446 1177
rect 1641 1172 1726 1177
rect 1809 1172 1974 1177
rect 1985 1172 2014 1177
rect 2081 1177 2086 1182
rect 2569 1177 2574 1182
rect 2081 1172 2110 1177
rect 2273 1172 2486 1177
rect 2513 1172 2574 1177
rect 2729 1177 2734 1182
rect 2729 1172 2758 1177
rect 1417 1167 1422 1172
rect 153 1162 302 1167
rect 561 1162 822 1167
rect 841 1162 982 1167
rect 1281 1162 1422 1167
rect 1473 1162 1614 1167
rect 1801 1162 1854 1167
rect 1937 1162 2022 1167
rect 2033 1162 2078 1167
rect 2129 1162 2254 1167
rect 2329 1162 2438 1167
rect 2625 1162 2830 1167
rect 841 1157 846 1162
rect 393 1152 550 1157
rect 601 1152 846 1157
rect 977 1157 982 1162
rect 2129 1157 2134 1162
rect 977 1152 1038 1157
rect 1737 1152 2134 1157
rect 2249 1157 2254 1162
rect 2249 1152 2358 1157
rect 2497 1152 2838 1157
rect 2857 1152 3054 1157
rect 2857 1147 2862 1152
rect 681 1142 966 1147
rect 1049 1142 1254 1147
rect 1289 1142 1454 1147
rect 497 1137 630 1142
rect 961 1137 1054 1142
rect 0 1132 502 1137
rect 625 1132 726 1137
rect 721 1127 726 1132
rect 825 1132 870 1137
rect 825 1127 830 1132
rect 1289 1127 1294 1142
rect 1449 1127 1454 1142
rect 1521 1142 1718 1147
rect 2017 1142 2070 1147
rect 2145 1142 2286 1147
rect 2297 1142 2366 1147
rect 2385 1142 2478 1147
rect 2497 1142 2630 1147
rect 2673 1142 2702 1147
rect 2833 1142 2862 1147
rect 3049 1147 3054 1152
rect 3049 1142 3080 1147
rect 1521 1137 1526 1142
rect 1713 1137 1894 1142
rect 2385 1137 2390 1142
rect 1497 1132 1526 1137
rect 1889 1132 1990 1137
rect 2129 1132 2174 1137
rect 2233 1132 2390 1137
rect 2473 1137 2478 1142
rect 2697 1137 2838 1142
rect 2473 1132 2662 1137
rect 2169 1127 2174 1132
rect 513 1122 614 1127
rect 721 1122 830 1127
rect 849 1122 942 1127
rect 961 1122 1214 1127
rect 1265 1122 1294 1127
rect 1313 1122 1382 1127
rect 1449 1122 1878 1127
rect 2113 1122 2166 1127
rect 2169 1122 3080 1127
rect 1313 1117 1318 1122
rect 1241 1112 1318 1117
rect 1377 1117 1382 1122
rect 1873 1117 1990 1122
rect 2113 1117 2118 1122
rect 1377 1112 1406 1117
rect 1441 1112 1566 1117
rect 1985 1112 2118 1117
rect 2161 1117 2166 1122
rect 2161 1112 2230 1117
rect 2273 1112 2406 1117
rect 2553 1112 2598 1117
rect 1585 1107 1718 1112
rect 2273 1107 2278 1112
rect 2401 1107 2558 1112
rect 265 1102 702 1107
rect 1089 1102 1174 1107
rect 1193 1102 1358 1107
rect 1457 1102 1590 1107
rect 1713 1102 1742 1107
rect 1761 1102 1910 1107
rect 2137 1102 2278 1107
rect 2289 1102 2366 1107
rect 2577 1102 2606 1107
rect 1089 1097 1094 1102
rect 721 1092 910 1097
rect 1065 1092 1094 1097
rect 1169 1097 1174 1102
rect 1353 1097 1462 1102
rect 1761 1097 1766 1102
rect 1169 1092 1334 1097
rect 721 1087 726 1092
rect 681 1082 726 1087
rect 905 1087 910 1092
rect 1329 1087 1334 1092
rect 1481 1092 1766 1097
rect 1905 1097 1910 1102
rect 2601 1097 2606 1102
rect 2801 1102 3080 1107
rect 2801 1097 2806 1102
rect 1905 1092 1966 1097
rect 2409 1092 2550 1097
rect 2601 1092 2806 1097
rect 1481 1087 1486 1092
rect 905 1082 1206 1087
rect 1329 1082 1486 1087
rect 1505 1082 1894 1087
rect 1889 1077 1894 1082
rect 1977 1082 2126 1087
rect 1977 1077 1982 1082
rect 0 1072 894 1077
rect 1201 1072 1230 1077
rect 1225 1067 1230 1072
rect 1577 1072 1742 1077
rect 1577 1067 1582 1072
rect 1737 1067 1742 1072
rect 1841 1072 1870 1077
rect 1889 1072 1982 1077
rect 2121 1077 2126 1082
rect 2185 1082 2214 1087
rect 2825 1082 2854 1087
rect 2185 1077 2190 1082
rect 2121 1072 2190 1077
rect 1841 1067 1846 1072
rect 1225 1062 1582 1067
rect 1601 1062 1630 1067
rect 1625 1057 1630 1062
rect 1689 1062 1718 1067
rect 1737 1062 1846 1067
rect 2209 1067 2214 1082
rect 2849 1077 2854 1082
rect 3049 1082 3080 1087
rect 3049 1077 3054 1082
rect 2297 1072 2446 1077
rect 2465 1072 2542 1077
rect 2849 1072 3054 1077
rect 2209 1062 2302 1067
rect 1689 1057 1694 1062
rect 1625 1052 1694 1057
rect 2209 1052 2246 1057
rect 2265 1047 2350 1052
rect 1809 1042 1950 1047
rect 1809 1037 1814 1042
rect 529 1032 566 1037
rect 585 1032 694 1037
rect 1449 1032 1718 1037
rect 1785 1032 1814 1037
rect 1945 1037 1950 1042
rect 1985 1042 2190 1047
rect 2217 1042 2270 1047
rect 2345 1042 2430 1047
rect 2617 1042 2678 1047
rect 2721 1042 2926 1047
rect 1985 1037 1990 1042
rect 1945 1032 1990 1037
rect 2185 1037 2190 1042
rect 2721 1037 2726 1042
rect 2185 1032 2334 1037
rect 481 1022 614 1027
rect 785 1017 790 1027
rect 889 1022 1022 1027
rect 1209 1022 1350 1027
rect 1209 1017 1214 1022
rect 0 1012 326 1017
rect 465 1012 790 1017
rect 1153 1012 1214 1017
rect 1345 1017 1350 1022
rect 1449 1017 1454 1032
rect 1345 1012 1374 1017
rect 1409 1007 1414 1017
rect 1425 1012 1454 1017
rect 1713 1017 1718 1032
rect 2329 1027 2334 1032
rect 2441 1032 2606 1037
rect 2441 1027 2446 1032
rect 1817 1022 1934 1027
rect 2081 1022 2174 1027
rect 2081 1017 2086 1022
rect 1713 1012 1774 1017
rect 2001 1012 2086 1017
rect 2169 1017 2174 1022
rect 2233 1022 2310 1027
rect 2329 1022 2446 1027
rect 2601 1027 2606 1032
rect 2689 1032 2726 1037
rect 2921 1037 2926 1042
rect 2921 1032 2950 1037
rect 3009 1032 3080 1037
rect 2689 1027 2694 1032
rect 2601 1022 2694 1027
rect 2737 1022 2806 1027
rect 2233 1017 2238 1022
rect 2169 1012 2238 1017
rect 2801 1017 2806 1022
rect 2801 1012 3080 1017
rect 1241 1002 1510 1007
rect 1609 1002 1702 1007
rect 2001 997 2006 1012
rect 2281 1002 2326 1007
rect 2417 1002 2582 1007
rect 393 992 542 997
rect 1225 992 1310 997
rect 1329 992 1462 997
rect 1473 992 1558 997
rect 1649 992 1830 997
rect 1889 992 2006 997
rect 2105 992 2270 997
rect 1457 987 1462 992
rect 1825 987 1830 992
rect 2265 987 2270 992
rect 2337 992 2486 997
rect 2569 992 2790 997
rect 2337 987 2342 992
rect 305 982 374 987
rect 305 977 310 982
rect 0 972 310 977
rect 369 977 374 982
rect 561 982 678 987
rect 929 982 1230 987
rect 561 977 566 982
rect 369 972 566 977
rect 673 977 678 982
rect 1225 977 1230 982
rect 1345 982 1414 987
rect 1457 982 1806 987
rect 1825 982 2030 987
rect 2265 982 2342 987
rect 2785 987 2790 992
rect 3049 992 3080 997
rect 3049 987 3054 992
rect 2785 982 3054 987
rect 1345 977 1350 982
rect 673 972 702 977
rect 1225 972 1350 977
rect 1393 972 1526 977
rect 1705 972 2038 977
rect 1081 962 1110 967
rect 1105 957 1110 962
rect 1177 962 1206 967
rect 1417 962 1782 967
rect 1945 962 1974 967
rect 2697 962 2766 967
rect 1177 957 1182 962
rect 1777 957 1950 962
rect 321 952 670 957
rect 777 952 870 957
rect 897 952 1014 957
rect 1105 952 1182 957
rect 1369 952 1470 957
rect 1665 952 1758 957
rect 641 942 758 947
rect 1513 942 1654 947
rect 1769 942 2022 947
rect 2361 942 2470 947
rect 2649 942 2678 947
rect 753 937 758 942
rect 1649 937 1774 942
rect 393 932 462 937
rect 753 932 942 937
rect 2241 932 2342 937
rect 2241 927 2246 932
rect 25 922 374 927
rect 25 917 30 922
rect 0 912 30 917
rect 369 917 374 922
rect 481 922 622 927
rect 953 922 1094 927
rect 1113 922 1270 927
rect 1337 922 1494 927
rect 1561 922 1734 927
rect 481 917 486 922
rect 369 912 486 917
rect 617 917 622 922
rect 1089 917 1094 922
rect 1337 917 1342 922
rect 617 912 822 917
rect 1089 912 1110 917
rect 1105 907 1110 912
rect 1281 912 1342 917
rect 1489 917 1494 922
rect 1729 917 1734 922
rect 1865 922 1894 927
rect 2225 922 2246 927
rect 2337 927 2342 932
rect 2337 922 3080 927
rect 1865 917 1870 922
rect 1489 912 1606 917
rect 1729 912 1870 917
rect 1961 912 2054 917
rect 2225 912 2230 922
rect 1281 907 1286 912
rect 1601 907 1606 912
rect 1001 902 1078 907
rect 1105 902 1286 907
rect 1353 902 1502 907
rect 1601 902 1638 907
rect 2025 902 2518 907
rect 0 892 622 897
rect 1073 887 1078 902
rect 1353 887 1358 902
rect 1497 897 1590 902
rect 2513 897 2518 902
rect 2745 902 2774 907
rect 2937 902 2966 907
rect 2745 897 2750 902
rect 1585 892 1710 897
rect 2513 892 2750 897
rect 2961 897 2966 902
rect 3049 902 3080 907
rect 3049 897 3054 902
rect 2961 892 3054 897
rect 1073 882 1358 887
rect 1377 882 1462 887
rect 1497 882 1574 887
rect 1569 877 1574 882
rect 1721 882 1782 887
rect 1721 877 1726 882
rect 0 872 446 877
rect 441 867 446 872
rect 601 872 630 877
rect 1569 872 1726 877
rect 2017 872 2094 877
rect 2241 872 2494 877
rect 601 867 606 872
rect 441 862 606 867
rect 945 862 1022 867
rect 2513 862 2686 867
rect 2241 857 2406 862
rect 2513 857 2518 862
rect 0 852 30 857
rect 25 847 30 852
rect 393 852 422 857
rect 1321 852 1630 857
rect 2217 852 2246 857
rect 2401 852 2430 857
rect 2441 852 2518 857
rect 2681 857 2686 862
rect 2681 852 2966 857
rect 393 847 398 852
rect 25 842 398 847
rect 1057 842 1318 847
rect 1633 842 1742 847
rect 1761 842 2454 847
rect 1313 837 1430 842
rect 1425 832 1454 837
rect 2313 832 2382 837
rect 2465 832 2670 837
rect 2377 827 2470 832
rect 1377 822 1414 827
rect 2057 822 2230 827
rect 2745 822 2838 827
rect 1377 817 1382 822
rect 0 812 318 817
rect 1177 812 1382 817
rect 2225 817 2230 822
rect 2225 812 2702 817
rect 2841 812 2870 817
rect 2937 812 3080 817
rect 2721 807 2846 812
rect 1025 802 1126 807
rect 1169 802 1238 807
rect 2169 802 2230 807
rect 2305 802 2382 807
rect 2657 802 2726 807
rect 353 792 942 797
rect 1513 792 1558 797
rect 2057 792 2166 797
rect 2225 792 2230 802
rect 2401 797 2526 802
rect 2657 797 2662 802
rect 2353 792 2406 797
rect 2521 792 2662 797
rect 2673 792 2982 797
rect 2161 787 2166 792
rect 1081 782 1214 787
rect 1257 782 1374 787
rect 1257 777 1262 782
rect 1097 772 1206 777
rect 1233 772 1262 777
rect 1369 777 1374 782
rect 1577 782 1646 787
rect 1737 782 1814 787
rect 2161 782 2510 787
rect 1577 777 1582 782
rect 1369 772 1398 777
rect 1433 772 1582 777
rect 1641 777 1646 782
rect 1641 772 1806 777
rect 425 762 494 767
rect 2017 762 2142 767
rect 425 757 430 762
rect 401 752 430 757
rect 489 757 494 762
rect 1297 757 1614 762
rect 2017 757 2022 762
rect 489 752 646 757
rect 889 752 918 757
rect 1137 752 1166 757
rect 1161 747 1166 752
rect 1273 752 1302 757
rect 1609 752 1886 757
rect 1953 752 2022 757
rect 2137 757 2142 762
rect 2137 752 2214 757
rect 2305 752 2358 757
rect 2577 752 2582 792
rect 2977 787 2982 792
rect 3049 792 3080 797
rect 3049 787 3054 792
rect 2977 782 3054 787
rect 2769 772 2958 777
rect 1273 747 1278 752
rect 2305 747 2310 752
rect 257 742 534 747
rect 529 727 534 742
rect 657 742 742 747
rect 969 742 1014 747
rect 1161 742 1278 747
rect 1329 742 1414 747
rect 1473 742 1526 747
rect 1569 742 1598 747
rect 657 727 662 742
rect 1329 737 1334 742
rect 1593 737 1702 742
rect 1833 737 1838 747
rect 1961 742 2054 747
rect 2065 742 2310 747
rect 2329 742 2382 747
rect 2473 742 2542 747
rect 2673 742 2918 747
rect 841 732 878 737
rect 153 722 246 727
rect 241 717 246 722
rect 353 722 510 727
rect 529 722 662 727
rect 873 727 878 732
rect 937 732 966 737
rect 1017 732 1110 737
rect 1297 732 1334 737
rect 1697 732 1950 737
rect 937 727 942 732
rect 1945 727 1950 732
rect 2065 727 2070 742
rect 2937 732 3054 737
rect 2625 727 2726 732
rect 2937 727 2942 732
rect 873 722 942 727
rect 1633 722 1662 727
rect 1945 722 2070 727
rect 2425 722 2630 727
rect 2721 722 2942 727
rect 3049 727 3054 732
rect 3049 722 3080 727
rect 353 717 358 722
rect 1633 717 1638 722
rect 241 712 358 717
rect 1153 712 1334 717
rect 1377 712 1454 717
rect 1609 712 1638 717
rect 1697 712 1822 717
rect 2225 712 2294 717
rect 1489 707 1574 712
rect 2225 707 2230 712
rect 377 702 470 707
rect 1417 702 1494 707
rect 1569 702 1598 707
rect 1593 697 1598 702
rect 1785 702 2230 707
rect 2289 707 2294 712
rect 2641 712 2710 717
rect 2289 702 2414 707
rect 1785 697 1790 702
rect 2409 697 2414 702
rect 2641 697 2646 712
rect 2705 707 2710 712
rect 2953 712 2990 717
rect 2953 707 2958 712
rect 2657 702 2686 707
rect 2705 702 2958 707
rect 3001 702 3080 707
rect 545 692 766 697
rect 905 692 942 697
rect 1385 692 1414 697
rect 1505 692 1534 697
rect 1593 692 1790 697
rect 1809 692 1838 697
rect 2409 692 2646 697
rect 1529 677 1534 692
rect 1809 677 1814 692
rect 2681 687 2686 702
rect 3001 687 3006 702
rect 2241 682 2278 687
rect 2681 682 3006 687
rect 1529 672 1814 677
rect 2153 672 2230 677
rect 1265 652 1438 657
rect 1265 647 1270 652
rect 273 642 446 647
rect 457 642 614 647
rect 945 642 1270 647
rect 1417 642 1902 647
rect 2641 642 2766 647
rect 2641 637 2646 642
rect 1393 632 1486 637
rect 2585 632 2646 637
rect 2761 637 2766 642
rect 2761 632 2790 637
rect 209 622 262 627
rect 257 617 262 622
rect 625 622 934 627
rect 625 617 630 622
rect 257 612 630 617
rect 929 617 934 622
rect 1281 622 1414 627
rect 1505 622 1550 627
rect 1921 622 1982 627
rect 2737 622 2758 627
rect 2969 622 3054 627
rect 1281 617 1286 622
rect 929 612 1286 617
rect 1409 617 1414 622
rect 2969 617 2974 622
rect 1409 612 1806 617
rect 1817 612 1902 617
rect 1969 612 2334 617
rect 2657 612 2686 617
rect 1969 607 1974 612
rect 1305 602 1446 607
rect 1769 602 1974 607
rect 2681 607 2686 612
rect 2801 612 2974 617
rect 3049 617 3054 622
rect 3049 612 3080 617
rect 2801 607 2806 612
rect 2681 602 2806 607
rect 657 592 766 597
rect 785 592 886 597
rect 1441 592 1446 602
rect 1545 597 1646 602
rect 1521 592 1550 597
rect 1641 592 1670 597
rect 1777 592 1862 597
rect 2017 592 2126 597
rect 2985 592 3080 597
rect 657 587 662 592
rect 305 582 614 587
rect 633 582 662 587
rect 761 587 766 592
rect 761 582 878 587
rect 1249 582 1334 587
rect 1465 582 1758 587
rect 609 577 614 582
rect 1753 577 1758 582
rect 1873 582 2078 587
rect 2225 582 2326 587
rect 1873 577 1878 582
rect 2225 577 2230 582
rect 609 572 630 577
rect 625 567 630 572
rect 745 572 798 577
rect 745 567 750 572
rect 625 562 750 567
rect 793 567 798 572
rect 897 572 1262 577
rect 1753 572 1878 577
rect 2201 572 2230 577
rect 2321 577 2326 582
rect 2321 572 2534 577
rect 897 567 902 572
rect 1561 567 1662 572
rect 1977 567 2062 572
rect 2529 567 2534 572
rect 793 562 902 567
rect 1201 562 1358 567
rect 1409 562 1566 567
rect 1657 562 1686 567
rect 1953 562 1982 567
rect 2057 562 2190 567
rect 2529 562 2822 567
rect 1953 557 1958 562
rect 2185 557 2278 562
rect 1577 552 1702 557
rect 1897 552 1958 557
rect 1977 552 2046 557
rect 2273 552 2358 557
rect 289 542 366 547
rect 553 542 606 547
rect 1041 542 1070 547
rect 1313 542 1438 547
rect 1497 542 1582 547
rect 289 537 294 542
rect 265 532 294 537
rect 361 537 366 542
rect 1577 537 1582 542
rect 1681 542 1710 547
rect 1769 542 1894 547
rect 2089 542 2222 547
rect 2273 542 2278 552
rect 2353 547 2358 552
rect 2385 552 2462 557
rect 2385 547 2390 552
rect 2289 542 2342 547
rect 2353 542 2390 547
rect 2401 542 2574 547
rect 2657 542 2838 547
rect 2865 542 2942 547
rect 1681 537 1686 542
rect 2833 537 2838 542
rect 361 532 390 537
rect 1201 532 1294 537
rect 1505 532 1558 537
rect 1577 532 1686 537
rect 1761 532 1790 537
rect 1905 532 2134 537
rect 1201 527 1206 532
rect 1177 522 1206 527
rect 1289 527 1294 532
rect 1785 527 1910 532
rect 2129 527 2134 532
rect 2585 532 2822 537
rect 2833 532 2862 537
rect 1289 522 1342 527
rect 1377 522 1486 527
rect 2129 522 2382 527
rect 1377 517 1382 522
rect 65 512 1278 517
rect 1273 507 1278 512
rect 1353 512 1382 517
rect 1481 517 1486 522
rect 2377 517 2382 522
rect 2585 517 2590 532
rect 2873 522 2990 527
rect 1481 512 2110 517
rect 2377 512 2590 517
rect 2657 512 2694 517
rect 1353 507 1358 512
rect 1273 502 1358 507
rect 1393 502 1494 507
rect 2257 502 2358 507
rect 2761 502 2862 507
rect 289 482 2046 487
rect 2513 482 2742 487
rect 2513 467 2518 482
rect 961 462 1062 467
rect 1641 462 1694 467
rect 2489 462 2518 467
rect 2737 467 2742 482
rect 2737 462 2782 467
rect 433 452 654 457
rect 1465 452 1622 457
rect 313 442 414 447
rect 313 437 318 442
rect 65 432 318 437
rect 409 437 414 442
rect 1353 442 1422 447
rect 1353 437 1358 442
rect 409 432 486 437
rect 1329 432 1358 437
rect 1417 437 1422 442
rect 1465 437 1470 452
rect 1617 447 1622 452
rect 1929 452 2758 457
rect 1929 447 1934 452
rect 1617 442 1702 447
rect 1697 437 1702 442
rect 1713 442 1934 447
rect 1713 437 1718 442
rect 2569 437 2654 442
rect 1417 432 1470 437
rect 1513 432 1598 437
rect 1697 432 1718 437
rect 1873 432 2046 437
rect 2257 432 2374 437
rect 2449 432 2574 437
rect 2649 432 2678 437
rect 2721 432 2766 437
rect 2857 432 2950 437
rect 1513 427 1518 432
rect 1409 422 1518 427
rect 1593 427 1598 432
rect 2257 427 2262 432
rect 1593 422 1694 427
rect 1793 422 1990 427
rect 2057 422 2262 427
rect 2369 427 2374 432
rect 2857 427 2862 432
rect 2369 422 2390 427
rect 2401 422 2502 427
rect 2585 422 2614 427
rect 2777 422 2862 427
rect 2945 427 2950 432
rect 2945 422 2998 427
rect 1985 417 2062 422
rect 233 412 262 417
rect 257 407 262 412
rect 329 412 518 417
rect 985 412 1086 417
rect 1169 412 1206 417
rect 1265 412 1966 417
rect 2273 412 2366 417
rect 2385 412 2390 422
rect 2609 417 2782 422
rect 329 407 334 412
rect 257 402 334 407
rect 513 397 518 412
rect 1169 407 1174 412
rect 561 402 678 407
rect 1057 402 1174 407
rect 1193 402 1254 407
rect 1449 402 2494 407
rect 2665 402 2694 407
rect 561 397 566 402
rect 513 392 566 397
rect 673 397 678 402
rect 1249 397 1454 402
rect 2689 397 2694 402
rect 2785 402 2934 407
rect 2785 397 2790 402
rect 673 392 806 397
rect 1049 392 1102 397
rect 1129 392 1230 397
rect 1473 392 1662 397
rect 1681 392 1750 397
rect 2297 392 2486 397
rect 2537 392 2646 397
rect 2689 392 2790 397
rect 1769 387 1902 392
rect 353 382 510 387
rect 729 382 782 387
rect 1201 382 1774 387
rect 1897 382 2342 387
rect 729 377 734 382
rect 2337 377 2342 382
rect 2569 382 2598 387
rect 2809 382 2926 387
rect 2569 377 2574 382
rect 577 372 734 377
rect 761 372 894 377
rect 1425 372 1446 377
rect 1569 372 1606 377
rect 1665 372 1734 377
rect 1785 372 1862 377
rect 2089 372 2230 377
rect 2337 372 2574 377
rect 577 367 582 372
rect 305 362 374 367
rect 433 362 582 367
rect 1209 362 1310 367
rect 1657 362 1718 367
rect 1905 362 2110 367
rect 433 337 438 362
rect 1209 357 1214 362
rect 753 352 894 357
rect 1185 352 1214 357
rect 1305 357 1310 362
rect 1305 352 1678 357
rect 1705 352 1726 357
rect 1777 352 1950 357
rect 1969 352 2086 357
rect 2121 352 2150 357
rect 2161 352 2590 357
rect 2161 347 2166 352
rect 505 342 678 347
rect 689 342 782 347
rect 969 342 1014 347
rect 1209 342 1294 347
rect 1497 342 1542 347
rect 1593 342 1654 347
rect 1961 342 1990 347
rect 2089 342 2166 347
rect 2865 342 2942 347
rect 217 332 438 337
rect 457 332 526 337
rect 673 327 678 342
rect 1985 337 2094 342
rect 761 332 790 337
rect 1409 332 1598 337
rect 1689 332 1918 337
rect 761 327 766 332
rect 1745 327 1750 332
rect 673 322 766 327
rect 1505 322 1566 327
rect 1673 322 1734 327
rect 1745 322 1782 327
rect 2025 322 2126 327
rect 2249 322 2310 327
rect 313 312 550 317
rect 1041 312 1078 317
rect 1785 312 1934 317
rect 2217 312 2278 317
rect 2385 312 2438 317
rect 2873 312 2998 317
rect 409 292 446 297
rect 489 292 782 297
rect 1609 292 1814 297
rect 1865 292 1910 297
rect 1921 292 1998 297
rect 2185 292 2374 297
rect 2385 292 2670 297
rect 1937 272 2270 277
rect 1201 252 1294 257
rect 1401 252 1574 257
rect 2137 252 2166 257
rect 1201 247 1206 252
rect 1041 242 1206 247
rect 1289 247 1294 252
rect 1289 242 1318 247
rect 393 232 518 237
rect 2033 232 2134 237
rect 1105 222 1134 227
rect 1209 222 1334 227
rect 1833 222 1902 227
rect 2089 222 2214 227
rect 2233 222 2358 227
rect 2401 222 2526 227
rect 2689 222 2806 227
rect 1833 217 1838 222
rect 1809 212 1838 217
rect 1897 217 1902 222
rect 1897 212 1926 217
rect 2881 212 2918 217
rect 2985 212 3080 217
rect 993 202 1038 207
rect 1369 202 1478 207
rect 1513 202 1614 207
rect 2881 197 2886 212
rect 1065 192 1414 197
rect 1505 192 1878 197
rect 1409 187 1510 192
rect 1873 187 1878 192
rect 1937 192 2886 197
rect 2897 192 2942 197
rect 1937 187 1942 192
rect 545 182 782 187
rect 1873 182 1942 187
rect 1369 172 1478 177
rect 1497 172 1550 177
rect 1697 172 1822 177
rect 2225 172 2278 177
rect 1209 162 1326 167
rect 1209 157 1214 162
rect 417 152 534 157
rect 833 152 894 157
rect 1185 152 1214 157
rect 1321 157 1326 162
rect 1369 157 1374 172
rect 1321 152 1374 157
rect 1473 157 1478 172
rect 1569 162 1654 167
rect 1569 157 1574 162
rect 1473 152 1574 157
rect 1649 157 1654 162
rect 1697 157 1702 172
rect 1649 152 1702 157
rect 1817 157 1822 172
rect 2113 162 2198 167
rect 2113 157 2118 162
rect 1817 152 2118 157
rect 2193 157 2198 162
rect 2417 162 2550 167
rect 2417 157 2422 162
rect 2193 152 2422 157
rect 2545 157 2550 162
rect 2593 162 2710 167
rect 2593 157 2598 162
rect 2545 152 2598 157
rect 2705 157 2710 162
rect 2753 162 2822 167
rect 2753 157 2758 162
rect 2705 152 2758 157
rect 2817 157 2822 162
rect 2817 152 2846 157
rect 2865 152 2918 157
rect 417 137 422 152
rect 529 147 534 152
rect 529 142 862 147
rect 953 137 958 147
rect 1105 142 1158 147
rect 1201 142 1278 147
rect 329 132 422 137
rect 441 132 518 137
rect 513 127 518 132
rect 593 132 622 137
rect 737 132 830 137
rect 953 132 1094 137
rect 593 127 598 132
rect 513 122 598 127
rect 1089 127 1094 132
rect 1201 127 1206 142
rect 1273 137 1278 142
rect 1401 142 1494 147
rect 1505 142 1510 152
rect 1521 142 1774 147
rect 1401 137 1406 142
rect 1273 132 1406 137
rect 1489 137 1494 142
rect 1521 137 1526 142
rect 1769 137 1774 142
rect 1873 142 1902 147
rect 2129 142 2158 147
rect 1873 137 1878 142
rect 1489 132 1526 137
rect 1633 132 1670 137
rect 1769 132 1878 137
rect 2153 137 2158 142
rect 2281 142 2510 147
rect 2281 137 2286 142
rect 2153 132 2286 137
rect 2505 137 2510 142
rect 2601 142 2654 147
rect 2601 137 2606 142
rect 2505 132 2606 137
rect 2649 137 2654 142
rect 2737 142 2790 147
rect 2737 137 2742 142
rect 2649 132 2742 137
rect 2785 137 2790 142
rect 2865 137 2870 152
rect 2897 142 2942 147
rect 2785 132 2870 137
rect 1089 122 1206 127
rect 1585 122 1614 127
rect 1681 122 1750 127
rect 2985 122 3080 127
rect 977 112 1022 117
rect 1793 112 1846 117
rect 321 102 590 107
rect 665 102 894 107
rect 569 92 678 97
rect 1465 92 1606 97
rect 361 82 630 87
rect 257 72 406 77
rect 401 67 406 72
rect 481 72 534 77
rect 481 67 486 72
rect 401 62 486 67
rect 529 67 534 72
rect 633 72 774 77
rect 2249 72 2342 77
rect 633 67 638 72
rect 529 62 638 67
rect 1113 52 1158 57
rect 2953 22 3038 27
rect 137 12 166 17
rect 161 7 166 12
rect 1329 12 1670 17
rect 1329 7 1334 12
rect 161 2 1334 7
use AND2X2  AND2X2_0
timestamp 1714281807
transform 1 0 2352 0 1 2170
box -8 -3 40 105
use AND2X2  AND2X2_1
timestamp 1714281807
transform 1 0 1792 0 1 370
box -8 -3 40 105
use AND2X2  AND2X2_2
timestamp 1714281807
transform 1 0 2344 0 1 370
box -8 -3 40 105
use AND2X2  AND2X2_3
timestamp 1714281807
transform 1 0 1928 0 1 370
box -8 -3 40 105
use AND2X2  AND2X2_4
timestamp 1714281807
transform 1 0 1464 0 1 370
box -8 -3 40 105
use AND2X2  AND2X2_5
timestamp 1714281807
transform 1 0 1200 0 1 370
box -8 -3 40 105
use AND2X2  AND2X2_6
timestamp 1714281807
transform 1 0 1208 0 -1 970
box -8 -3 40 105
use AND2X2  AND2X2_7
timestamp 1714281807
transform 1 0 1744 0 1 1170
box -8 -3 40 105
use AND2X2  AND2X2_8
timestamp 1714281807
transform 1 0 1672 0 1 1570
box -8 -3 40 105
use AND2X2  AND2X2_9
timestamp 1714281807
transform 1 0 936 0 1 1370
box -8 -3 40 105
use AND2X2  AND2X2_10
timestamp 1714281807
transform 1 0 2224 0 1 1770
box -8 -3 40 105
use AND2X2  AND2X2_11
timestamp 1714281807
transform 1 0 2680 0 1 1970
box -8 -3 40 105
use AND2X2  AND2X2_12
timestamp 1714281807
transform 1 0 2216 0 1 2570
box -8 -3 40 105
use AND2X2  AND2X2_13
timestamp 1714281807
transform 1 0 1640 0 1 2570
box -8 -3 40 105
use AND2X2  AND2X2_14
timestamp 1714281807
transform 1 0 984 0 -1 1770
box -8 -3 40 105
use AND2X2  AND2X2_15
timestamp 1714281807
transform 1 0 2568 0 1 2570
box -8 -3 40 105
use AND2X2  AND2X2_16
timestamp 1714281807
transform 1 0 1352 0 1 2570
box -8 -3 40 105
use AND2X2  AND2X2_17
timestamp 1714281807
transform 1 0 2544 0 1 1170
box -8 -3 40 105
use AND2X2  AND2X2_18
timestamp 1714281807
transform 1 0 2192 0 1 1170
box -8 -3 40 105
use AND2X2  AND2X2_19
timestamp 1714281807
transform 1 0 992 0 1 1370
box -8 -3 40 105
use AND2X2  AND2X2_20
timestamp 1714281807
transform 1 0 864 0 -1 1370
box -8 -3 40 105
use AND2X2  AND2X2_21
timestamp 1714281807
transform 1 0 2608 0 -1 570
box -8 -3 40 105
use AND2X2  AND2X2_22
timestamp 1714281807
transform 1 0 968 0 -1 1370
box -8 -3 40 105
use AND2X2  AND2X2_23
timestamp 1714281807
transform 1 0 896 0 -1 1370
box -8 -3 40 105
use AND2X2  AND2X2_24
timestamp 1714281807
transform 1 0 1832 0 1 1970
box -8 -3 40 105
use AND2X2  AND2X2_25
timestamp 1714281807
transform 1 0 848 0 -1 770
box -8 -3 40 105
use AOI21X1  AOI21X1_0
timestamp 1714281807
transform 1 0 776 0 -1 2770
box -7 -3 39 105
use AOI21X1  AOI21X1_1
timestamp 1714281807
transform 1 0 608 0 -1 2770
box -7 -3 39 105
use AOI21X1  AOI21X1_2
timestamp 1714281807
transform 1 0 408 0 1 2770
box -7 -3 39 105
use AOI21X1  AOI21X1_3
timestamp 1714281807
transform 1 0 496 0 -1 2970
box -7 -3 39 105
use AOI21X1  AOI21X1_4
timestamp 1714281807
transform 1 0 696 0 -1 2970
box -7 -3 39 105
use AOI21X1  AOI21X1_5
timestamp 1714281807
transform 1 0 856 0 -1 2970
box -7 -3 39 105
use AOI21X1  AOI21X1_6
timestamp 1714281807
transform 1 0 432 0 -1 570
box -7 -3 39 105
use AOI21X1  AOI21X1_7
timestamp 1714281807
transform 1 0 400 0 -1 370
box -7 -3 39 105
use AOI21X1  AOI21X1_8
timestamp 1714281807
transform 1 0 744 0 1 170
box -7 -3 39 105
use AOI21X1  AOI21X1_9
timestamp 1714281807
transform 1 0 800 0 -1 170
box -7 -3 39 105
use AOI22X1  AOI22X1_0
timestamp 1714281807
transform 1 0 2456 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_1
timestamp 1714281807
transform 1 0 2528 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_2
timestamp 1714281807
transform 1 0 2264 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_3
timestamp 1714281807
transform 1 0 1120 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_4
timestamp 1714281807
transform 1 0 1992 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_5
timestamp 1714281807
transform 1 0 2080 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_6
timestamp 1714281807
transform 1 0 1872 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_7
timestamp 1714281807
transform 1 0 1088 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_8
timestamp 1714281807
transform 1 0 1528 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_9
timestamp 1714281807
transform 1 0 1688 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_10
timestamp 1714281807
transform 1 0 1408 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_11
timestamp 1714281807
transform 1 0 1144 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_12
timestamp 1714281807
transform 1 0 1128 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_13
timestamp 1714281807
transform 1 0 1176 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_14
timestamp 1714281807
transform 1 0 1264 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_15
timestamp 1714281807
transform 1 0 1016 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_16
timestamp 1714281807
transform 1 0 1176 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_17
timestamp 1714281807
transform 1 0 1168 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_18
timestamp 1714281807
transform 1 0 1224 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_19
timestamp 1714281807
transform 1 0 992 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_20
timestamp 1714281807
transform 1 0 1824 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_21
timestamp 1714281807
transform 1 0 1688 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_22
timestamp 1714281807
transform 1 0 1760 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_23
timestamp 1714281807
transform 1 0 1096 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_24
timestamp 1714281807
transform 1 0 1640 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_25
timestamp 1714281807
transform 1 0 1648 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_26
timestamp 1714281807
transform 1 0 1728 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_27
timestamp 1714281807
transform 1 0 1184 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_28
timestamp 1714281807
transform 1 0 2232 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_29
timestamp 1714281807
transform 1 0 2320 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_30
timestamp 1714281807
transform 1 0 2312 0 1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_31
timestamp 1714281807
transform 1 0 1264 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_32
timestamp 1714281807
transform 1 0 2744 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_33
timestamp 1714281807
transform 1 0 2720 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_34
timestamp 1714281807
transform 1 0 2800 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_35
timestamp 1714281807
transform 1 0 1352 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_36
timestamp 1714281807
transform 1 0 2280 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_37
timestamp 1714281807
transform 1 0 2096 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_38
timestamp 1714281807
transform 1 0 2368 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_39
timestamp 1714281807
transform 1 0 1360 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_40
timestamp 1714281807
transform 1 0 1792 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_41
timestamp 1714281807
transform 1 0 1712 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_42
timestamp 1714281807
transform 1 0 1912 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_43
timestamp 1714281807
transform 1 0 1272 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_44
timestamp 1714281807
transform 1 0 2696 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_45
timestamp 1714281807
transform 1 0 2504 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_46
timestamp 1714281807
transform 1 0 2784 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_47
timestamp 1714281807
transform 1 0 1264 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_48
timestamp 1714281807
transform 1 0 1408 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_49
timestamp 1714281807
transform 1 0 1456 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_50
timestamp 1714281807
transform 1 0 1384 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_51
timestamp 1714281807
transform 1 0 1272 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_52
timestamp 1714281807
transform 1 0 2736 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_53
timestamp 1714281807
transform 1 0 2544 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_54
timestamp 1714281807
transform 1 0 2736 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_55
timestamp 1714281807
transform 1 0 1352 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_56
timestamp 1714281807
transform 1 0 2280 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_57
timestamp 1714281807
transform 1 0 2192 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_58
timestamp 1714281807
transform 1 0 2280 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_59
timestamp 1714281807
transform 1 0 1272 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_60
timestamp 1714281807
transform 1 0 2800 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_61
timestamp 1714281807
transform 1 0 2720 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_62
timestamp 1714281807
transform 1 0 2744 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_63
timestamp 1714281807
transform 1 0 1216 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_64
timestamp 1714281807
transform 1 0 776 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_65
timestamp 1714281807
transform 1 0 1928 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_66
timestamp 1714281807
transform 1 0 2008 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_67
timestamp 1714281807
transform 1 0 1936 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_68
timestamp 1714281807
transform 1 0 2032 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_69
timestamp 1714281807
transform 1 0 288 0 -1 370
box -8 -3 46 105
use BUFX2  BUFX2_0
timestamp 1714281807
transform 1 0 1000 0 -1 970
box -5 -3 28 105
use BUFX2  BUFX2_1
timestamp 1714281807
transform 1 0 2056 0 1 970
box -5 -3 28 105
use BUFX2  BUFX2_2
timestamp 1714281807
transform 1 0 1704 0 1 970
box -5 -3 28 105
use BUFX2  BUFX2_3
timestamp 1714281807
transform 1 0 1504 0 -1 970
box -5 -3 28 105
use BUFX2  BUFX2_4
timestamp 1714281807
transform 1 0 920 0 1 770
box -5 -3 28 105
use BUFX2  BUFX2_5
timestamp 1714281807
transform 1 0 2096 0 1 1770
box -5 -3 28 105
use BUFX2  BUFX2_6
timestamp 1714281807
transform 1 0 2136 0 -1 2370
box -5 -3 28 105
use BUFX2  BUFX2_7
timestamp 1714281807
transform 1 0 2080 0 1 970
box -5 -3 28 105
use BUFX2  BUFX2_8
timestamp 1714281807
transform 1 0 1728 0 1 970
box -5 -3 28 105
use BUFX2  BUFX2_9
timestamp 1714281807
transform 1 0 1728 0 1 1370
box -5 -3 28 105
use BUFX2  BUFX2_10
timestamp 1714281807
transform 1 0 1720 0 -1 1570
box -5 -3 28 105
use BUFX2  BUFX2_11
timestamp 1714281807
transform 1 0 1560 0 -1 970
box -5 -3 28 105
use BUFX2  BUFX2_12
timestamp 1714281807
transform 1 0 1528 0 -1 970
box -5 -3 28 105
use BUFX2  BUFX2_13
timestamp 1714281807
transform 1 0 1392 0 1 970
box -5 -3 28 105
use BUFX2  BUFX2_14
timestamp 1714281807
transform 1 0 944 0 1 770
box -5 -3 28 105
use BUFX2  BUFX2_15
timestamp 1714281807
transform 1 0 1232 0 1 1170
box -5 -3 28 105
use BUFX2  BUFX2_16
timestamp 1714281807
transform 1 0 1040 0 1 1170
box -5 -3 28 105
use BUFX2  BUFX2_17
timestamp 1714281807
transform 1 0 1208 0 1 1170
box -5 -3 28 105
use BUFX2  BUFX2_18
timestamp 1714281807
transform 1 0 1064 0 1 1170
box -5 -3 28 105
use BUFX2  BUFX2_19
timestamp 1714281807
transform 1 0 1240 0 -1 1370
box -5 -3 28 105
use BUFX2  BUFX2_20
timestamp 1714281807
transform 1 0 1272 0 -1 1370
box -5 -3 28 105
use BUFX2  BUFX2_21
timestamp 1714281807
transform 1 0 1376 0 -1 1370
box -5 -3 28 105
use BUFX2  BUFX2_22
timestamp 1714281807
transform 1 0 1344 0 -1 1370
box -5 -3 28 105
use BUFX2  BUFX2_23
timestamp 1714281807
transform 1 0 1320 0 -1 1370
box -5 -3 28 105
use BUFX2  BUFX2_24
timestamp 1714281807
transform 1 0 1016 0 -1 1170
box -5 -3 28 105
use BUFX2  BUFX2_25
timestamp 1714281807
transform 1 0 1184 0 1 1170
box -5 -3 28 105
use BUFX2  BUFX2_26
timestamp 1714281807
transform 1 0 2128 0 -1 1370
box -5 -3 28 105
use BUFX2  BUFX2_27
timestamp 1714281807
transform 1 0 2016 0 1 1370
box -5 -3 28 105
use BUFX2  BUFX2_28
timestamp 1714281807
transform 1 0 2112 0 -1 1570
box -5 -3 28 105
use BUFX2  BUFX2_29
timestamp 1714281807
transform 1 0 2152 0 -1 1370
box -5 -3 28 105
use DFFNEGX1  DFFNEGX1_0
timestamp 1714281807
transform 1 0 960 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_1
timestamp 1714281807
transform 1 0 1056 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_2
timestamp 1714281807
transform 1 0 744 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_3
timestamp 1714281807
transform 1 0 544 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_4
timestamp 1714281807
transform 1 0 320 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_5
timestamp 1714281807
transform 1 0 120 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_6
timestamp 1714281807
transform 1 0 96 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_7
timestamp 1714281807
transform 1 0 184 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_8
timestamp 1714281807
transform 1 0 360 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_9
timestamp 1714281807
transform 1 0 248 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_10
timestamp 1714281807
transform 1 0 432 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_11
timestamp 1714281807
transform 1 0 680 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_12
timestamp 1714281807
transform 1 0 840 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_13
timestamp 1714281807
transform 1 0 936 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_14
timestamp 1714281807
transform 1 0 688 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_15
timestamp 1714281807
transform 1 0 552 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_16
timestamp 1714281807
transform 1 0 592 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_17
timestamp 1714281807
transform 1 0 176 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_18
timestamp 1714281807
transform 1 0 152 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_19
timestamp 1714281807
transform 1 0 320 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_20
timestamp 1714281807
transform 1 0 816 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_21
timestamp 1714281807
transform 1 0 1008 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_22
timestamp 1714281807
transform 1 0 1160 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_23
timestamp 1714281807
transform 1 0 1216 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_24
timestamp 1714281807
transform 1 0 608 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_25
timestamp 1714281807
transform 1 0 592 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_26
timestamp 1714281807
transform 1 0 480 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_27
timestamp 1714281807
transform 1 0 504 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_28
timestamp 1714281807
transform 1 0 1104 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_29
timestamp 1714281807
transform 1 0 1064 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_30
timestamp 1714281807
transform 1 0 824 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_31
timestamp 1714281807
transform 1 0 960 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_32
timestamp 1714281807
transform 1 0 1176 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_33
timestamp 1714281807
transform 1 0 1200 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_34
timestamp 1714281807
transform 1 0 1288 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_35
timestamp 1714281807
transform 1 0 1296 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_36
timestamp 1714281807
transform 1 0 2584 0 1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_37
timestamp 1714281807
transform 1 0 2600 0 -1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_38
timestamp 1714281807
transform 1 0 2616 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_39
timestamp 1714281807
transform 1 0 1016 0 1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_40
timestamp 1714281807
transform 1 0 1048 0 -1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_41
timestamp 1714281807
transform 1 0 1088 0 1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_42
timestamp 1714281807
transform 1 0 1296 0 -1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_43
timestamp 1714281807
transform 1 0 824 0 1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_44
timestamp 1714281807
transform 1 0 688 0 1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_45
timestamp 1714281807
transform 1 0 1288 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_46
timestamp 1714281807
transform 1 0 784 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_47
timestamp 1714281807
transform 1 0 496 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_48
timestamp 1714281807
transform 1 0 264 0 -1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_49
timestamp 1714281807
transform 1 0 128 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_50
timestamp 1714281807
transform 1 0 96 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_51
timestamp 1714281807
transform 1 0 288 0 1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_52
timestamp 1714281807
transform 1 0 376 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_53
timestamp 1714281807
transform 1 0 312 0 -1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_54
timestamp 1714281807
transform 1 0 544 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_55
timestamp 1714281807
transform 1 0 2192 0 1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_56
timestamp 1714281807
transform 1 0 2112 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_57
timestamp 1714281807
transform 1 0 2392 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_58
timestamp 1714281807
transform 1 0 2664 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_59
timestamp 1714281807
transform 1 0 2760 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_60
timestamp 1714281807
transform 1 0 2640 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_61
timestamp 1714281807
transform 1 0 2072 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_62
timestamp 1714281807
transform 1 0 2168 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_63
timestamp 1714281807
transform 1 0 2296 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_64
timestamp 1714281807
transform 1 0 1744 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_65
timestamp 1714281807
transform 1 0 1832 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_66
timestamp 1714281807
transform 1 0 1848 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_67
timestamp 1714281807
transform 1 0 2488 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_68
timestamp 1714281807
transform 1 0 2680 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_69
timestamp 1714281807
transform 1 0 2600 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_70
timestamp 1714281807
transform 1 0 2432 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_71
timestamp 1714281807
transform 1 0 2568 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_72
timestamp 1714281807
transform 1 0 2664 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_73
timestamp 1714281807
transform 1 0 1904 0 -1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_74
timestamp 1714281807
transform 1 0 1960 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_75
timestamp 1714281807
transform 1 0 2016 0 -1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_76
timestamp 1714281807
transform 1 0 1888 0 -1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_77
timestamp 1714281807
transform 1 0 1936 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_78
timestamp 1714281807
transform 1 0 1880 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_79
timestamp 1714281807
transform 1 0 1416 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_80
timestamp 1714281807
transform 1 0 1240 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_81
timestamp 1714281807
transform 1 0 1312 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_82
timestamp 1714281807
transform 1 0 1472 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_83
timestamp 1714281807
transform 1 0 1432 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_84
timestamp 1714281807
transform 1 0 1392 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_85
timestamp 1714281807
transform 1 0 1248 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_86
timestamp 1714281807
transform 1 0 1584 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_87
timestamp 1714281807
transform 1 0 1256 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_88
timestamp 1714281807
transform 1 0 1800 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_89
timestamp 1714281807
transform 1 0 1888 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_90
timestamp 1714281807
transform 1 0 1728 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_91
timestamp 1714281807
transform 1 0 1800 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_92
timestamp 1714281807
transform 1 0 2136 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_93
timestamp 1714281807
transform 1 0 1920 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_94
timestamp 1714281807
transform 1 0 2264 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_95
timestamp 1714281807
transform 1 0 2448 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_96
timestamp 1714281807
transform 1 0 2376 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_97
timestamp 1714281807
transform 1 0 2344 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_98
timestamp 1714281807
transform 1 0 2304 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_99
timestamp 1714281807
transform 1 0 2384 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_100
timestamp 1714281807
transform 1 0 360 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_101
timestamp 1714281807
transform 1 0 360 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_102
timestamp 1714281807
transform 1 0 736 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_103
timestamp 1714281807
transform 1 0 536 0 -1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_104
timestamp 1714281807
transform 1 0 424 0 -1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_105
timestamp 1714281807
transform 1 0 312 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_106
timestamp 1714281807
transform 1 0 2424 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_107
timestamp 1714281807
transform 1 0 2408 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_108
timestamp 1714281807
transform 1 0 2336 0 -1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_109
timestamp 1714281807
transform 1 0 2904 0 1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_110
timestamp 1714281807
transform 1 0 2768 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_111
timestamp 1714281807
transform 1 0 2856 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_112
timestamp 1714281807
transform 1 0 2248 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_113
timestamp 1714281807
transform 1 0 2120 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_114
timestamp 1714281807
transform 1 0 2376 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_115
timestamp 1714281807
transform 1 0 2752 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_116
timestamp 1714281807
transform 1 0 2480 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_117
timestamp 1714281807
transform 1 0 2880 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_118
timestamp 1714281807
transform 1 0 1256 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_119
timestamp 1714281807
transform 1 0 1376 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_120
timestamp 1714281807
transform 1 0 1272 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_121
timestamp 1714281807
transform 1 0 2904 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_122
timestamp 1714281807
transform 1 0 2584 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_123
timestamp 1714281807
transform 1 0 2888 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_124
timestamp 1714281807
transform 1 0 2904 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_125
timestamp 1714281807
transform 1 0 2712 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_126
timestamp 1714281807
transform 1 0 2904 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_127
timestamp 1714281807
transform 1 0 2248 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_128
timestamp 1714281807
transform 1 0 2112 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_129
timestamp 1714281807
transform 1 0 2200 0 -1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_130
timestamp 1714281807
transform 1 0 1808 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_131
timestamp 1714281807
transform 1 0 1696 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_132
timestamp 1714281807
transform 1 0 1920 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_133
timestamp 1714281807
transform 1 0 1800 0 -1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_134
timestamp 1714281807
transform 1 0 1512 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_135
timestamp 1714281807
transform 1 0 1512 0 1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_136
timestamp 1714281807
transform 1 0 1864 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_137
timestamp 1714281807
transform 1 0 1576 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_138
timestamp 1714281807
transform 1 0 1840 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_139
timestamp 1714281807
transform 1 0 1272 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_140
timestamp 1714281807
transform 1 0 960 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_141
timestamp 1714281807
transform 1 0 968 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_142
timestamp 1714281807
transform 1 0 1240 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_143
timestamp 1714281807
transform 1 0 1056 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_144
timestamp 1714281807
transform 1 0 952 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_145
timestamp 1714281807
transform 1 0 1376 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_146
timestamp 1714281807
transform 1 0 1640 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_147
timestamp 1714281807
transform 1 0 1520 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_148
timestamp 1714281807
transform 1 0 1840 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_149
timestamp 1714281807
transform 1 0 1952 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_150
timestamp 1714281807
transform 1 0 2120 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_151
timestamp 1714281807
transform 1 0 2256 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_152
timestamp 1714281807
transform 1 0 2528 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_153
timestamp 1714281807
transform 1 0 2432 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_154
timestamp 1714281807
transform 1 0 1320 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_155
timestamp 1714281807
transform 1 0 920 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_156
timestamp 1714281807
transform 1 0 1856 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_157
timestamp 1714281807
transform 1 0 2168 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_158
timestamp 1714281807
transform 1 0 2168 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_159
timestamp 1714281807
transform 1 0 2064 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_160
timestamp 1714281807
transform 1 0 2080 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_161
timestamp 1714281807
transform 1 0 2024 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_162
timestamp 1714281807
transform 1 0 1512 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_163
timestamp 1714281807
transform 1 0 1464 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_164
timestamp 1714281807
transform 1 0 1520 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_165
timestamp 1714281807
transform 1 0 1512 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_166
timestamp 1714281807
transform 1 0 1656 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_167
timestamp 1714281807
transform 1 0 1520 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_168
timestamp 1714281807
transform 1 0 2008 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_169
timestamp 1714281807
transform 1 0 2072 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_170
timestamp 1714281807
transform 1 0 1560 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_171
timestamp 1714281807
transform 1 0 1824 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_172
timestamp 1714281807
transform 1 0 2160 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_173
timestamp 1714281807
transform 1 0 2176 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_174
timestamp 1714281807
transform 1 0 2344 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_175
timestamp 1714281807
transform 1 0 2568 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_176
timestamp 1714281807
transform 1 0 2576 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_177
timestamp 1714281807
transform 1 0 2776 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_178
timestamp 1714281807
transform 1 0 2856 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_179
timestamp 1714281807
transform 1 0 2848 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_180
timestamp 1714281807
transform 1 0 2112 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_181
timestamp 1714281807
transform 1 0 2536 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_182
timestamp 1714281807
transform 1 0 2280 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_183
timestamp 1714281807
transform 1 0 2528 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_184
timestamp 1714281807
transform 1 0 2872 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_185
timestamp 1714281807
transform 1 0 2776 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_186
timestamp 1714281807
transform 1 0 1616 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_187
timestamp 1714281807
transform 1 0 1648 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_188
timestamp 1714281807
transform 1 0 1608 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_189
timestamp 1714281807
transform 1 0 2464 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_190
timestamp 1714281807
transform 1 0 2816 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_191
timestamp 1714281807
transform 1 0 2872 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_192
timestamp 1714281807
transform 1 0 1744 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_193
timestamp 1714281807
transform 1 0 1992 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_194
timestamp 1714281807
transform 1 0 1976 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_195
timestamp 1714281807
transform 1 0 2072 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_196
timestamp 1714281807
transform 1 0 2232 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_197
timestamp 1714281807
transform 1 0 2344 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_198
timestamp 1714281807
transform 1 0 2864 0 1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_199
timestamp 1714281807
transform 1 0 2864 0 -1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_200
timestamp 1714281807
transform 1 0 2872 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_201
timestamp 1714281807
transform 1 0 2120 0 -1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_202
timestamp 1714281807
transform 1 0 1984 0 1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_203
timestamp 1714281807
transform 1 0 2144 0 1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_204
timestamp 1714281807
transform 1 0 1712 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_205
timestamp 1714281807
transform 1 0 1576 0 1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_206
timestamp 1714281807
transform 1 0 1608 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_207
timestamp 1714281807
transform 1 0 1744 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_208
timestamp 1714281807
transform 1 0 1624 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_209
timestamp 1714281807
transform 1 0 1728 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_210
timestamp 1714281807
transform 1 0 1064 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_211
timestamp 1714281807
transform 1 0 904 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_212
timestamp 1714281807
transform 1 0 912 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_213
timestamp 1714281807
transform 1 0 1056 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_214
timestamp 1714281807
transform 1 0 944 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_215
timestamp 1714281807
transform 1 0 912 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_216
timestamp 1714281807
transform 1 0 1240 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_217
timestamp 1714281807
transform 1 0 1576 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_218
timestamp 1714281807
transform 1 0 1416 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_219
timestamp 1714281807
transform 1 0 1736 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_220
timestamp 1714281807
transform 1 0 1888 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_221
timestamp 1714281807
transform 1 0 2120 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_222
timestamp 1714281807
transform 1 0 2296 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_223
timestamp 1714281807
transform 1 0 2616 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_224
timestamp 1714281807
transform 1 0 2472 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_225
timestamp 1714281807
transform 1 0 2752 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_226
timestamp 1714281807
transform 1 0 2904 0 -1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_227
timestamp 1714281807
transform 1 0 2904 0 1 170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_228
timestamp 1714281807
transform 1 0 2616 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_229
timestamp 1714281807
transform 1 0 2472 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_230
timestamp 1714281807
transform 1 0 2488 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_231
timestamp 1714281807
transform 1 0 2584 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_232
timestamp 1714281807
transform 1 0 2720 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_233
timestamp 1714281807
transform 1 0 2824 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_234
timestamp 1714281807
transform 1 0 1568 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_235
timestamp 1714281807
transform 1 0 1648 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_236
timestamp 1714281807
transform 1 0 1600 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_237
timestamp 1714281807
transform 1 0 2568 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_238
timestamp 1714281807
transform 1 0 2672 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_239
timestamp 1714281807
transform 1 0 2776 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_240
timestamp 1714281807
transform 1 0 1664 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_241
timestamp 1714281807
transform 1 0 1880 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_242
timestamp 1714281807
transform 1 0 1976 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_243
timestamp 1714281807
transform 1 0 2128 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_244
timestamp 1714281807
transform 1 0 2296 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_245
timestamp 1714281807
transform 1 0 2464 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_246
timestamp 1714281807
transform 1 0 2568 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_247
timestamp 1714281807
transform 1 0 2472 0 1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_248
timestamp 1714281807
transform 1 0 2512 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_249
timestamp 1714281807
transform 1 0 2480 0 -1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_250
timestamp 1714281807
transform 1 0 2480 0 1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_251
timestamp 1714281807
transform 1 0 2496 0 -1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_252
timestamp 1714281807
transform 1 0 1376 0 -1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_253
timestamp 1714281807
transform 1 0 1384 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_254
timestamp 1714281807
transform 1 0 1456 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_255
timestamp 1714281807
transform 1 0 1384 0 1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_256
timestamp 1714281807
transform 1 0 736 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_257
timestamp 1714281807
transform 1 0 712 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_258
timestamp 1714281807
transform 1 0 1416 0 -1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_259
timestamp 1714281807
transform 1 0 704 0 -1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_260
timestamp 1714281807
transform 1 0 88 0 1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_261
timestamp 1714281807
transform 1 0 120 0 -1 1570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_262
timestamp 1714281807
transform 1 0 216 0 -1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_263
timestamp 1714281807
transform 1 0 240 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_264
timestamp 1714281807
transform 1 0 152 0 1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_265
timestamp 1714281807
transform 1 0 200 0 -1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_266
timestamp 1714281807
transform 1 0 264 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_267
timestamp 1714281807
transform 1 0 232 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_268
timestamp 1714281807
transform 1 0 792 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_269
timestamp 1714281807
transform 1 0 296 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_270
timestamp 1714281807
transform 1 0 224 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_271
timestamp 1714281807
transform 1 0 352 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_272
timestamp 1714281807
transform 1 0 232 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_273
timestamp 1714281807
transform 1 0 560 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_274
timestamp 1714281807
transform 1 0 688 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_275
timestamp 1714281807
transform 1 0 760 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_276
timestamp 1714281807
transform 1 0 848 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_277
timestamp 1714281807
transform 1 0 824 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_278
timestamp 1714281807
transform 1 0 344 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_279
timestamp 1714281807
transform 1 0 536 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_280
timestamp 1714281807
transform 1 0 632 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_281
timestamp 1714281807
transform 1 0 440 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_282
timestamp 1714281807
transform 1 0 728 0 1 770
box -8 -3 104 105
use FILL  FILL_0
timestamp 1714281807
transform 1 0 3000 0 -1 2970
box -8 -3 16 105
use FILL  FILL_1
timestamp 1714281807
transform 1 0 2992 0 -1 2970
box -8 -3 16 105
use FILL  FILL_2
timestamp 1714281807
transform 1 0 2984 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3
timestamp 1714281807
transform 1 0 2976 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4
timestamp 1714281807
transform 1 0 2968 0 -1 2970
box -8 -3 16 105
use FILL  FILL_5
timestamp 1714281807
transform 1 0 2960 0 -1 2970
box -8 -3 16 105
use FILL  FILL_6
timestamp 1714281807
transform 1 0 2952 0 -1 2970
box -8 -3 16 105
use FILL  FILL_7
timestamp 1714281807
transform 1 0 2944 0 -1 2970
box -8 -3 16 105
use FILL  FILL_8
timestamp 1714281807
transform 1 0 2936 0 -1 2970
box -8 -3 16 105
use FILL  FILL_9
timestamp 1714281807
transform 1 0 2928 0 -1 2970
box -8 -3 16 105
use FILL  FILL_10
timestamp 1714281807
transform 1 0 2920 0 -1 2970
box -8 -3 16 105
use FILL  FILL_11
timestamp 1714281807
transform 1 0 2912 0 -1 2970
box -8 -3 16 105
use FILL  FILL_12
timestamp 1714281807
transform 1 0 2904 0 -1 2970
box -8 -3 16 105
use FILL  FILL_13
timestamp 1714281807
transform 1 0 2896 0 -1 2970
box -8 -3 16 105
use FILL  FILL_14
timestamp 1714281807
transform 1 0 2888 0 -1 2970
box -8 -3 16 105
use FILL  FILL_15
timestamp 1714281807
transform 1 0 2880 0 -1 2970
box -8 -3 16 105
use FILL  FILL_16
timestamp 1714281807
transform 1 0 2872 0 -1 2970
box -8 -3 16 105
use FILL  FILL_17
timestamp 1714281807
transform 1 0 2768 0 -1 2970
box -8 -3 16 105
use FILL  FILL_18
timestamp 1714281807
transform 1 0 2664 0 -1 2970
box -8 -3 16 105
use FILL  FILL_19
timestamp 1714281807
transform 1 0 2560 0 -1 2970
box -8 -3 16 105
use FILL  FILL_20
timestamp 1714281807
transform 1 0 2456 0 -1 2970
box -8 -3 16 105
use FILL  FILL_21
timestamp 1714281807
transform 1 0 2448 0 -1 2970
box -8 -3 16 105
use FILL  FILL_22
timestamp 1714281807
transform 1 0 2440 0 -1 2970
box -8 -3 16 105
use FILL  FILL_23
timestamp 1714281807
transform 1 0 2408 0 -1 2970
box -8 -3 16 105
use FILL  FILL_24
timestamp 1714281807
transform 1 0 2400 0 -1 2970
box -8 -3 16 105
use FILL  FILL_25
timestamp 1714281807
transform 1 0 2392 0 -1 2970
box -8 -3 16 105
use FILL  FILL_26
timestamp 1714281807
transform 1 0 2288 0 -1 2970
box -8 -3 16 105
use FILL  FILL_27
timestamp 1714281807
transform 1 0 2280 0 -1 2970
box -8 -3 16 105
use FILL  FILL_28
timestamp 1714281807
transform 1 0 2248 0 -1 2970
box -8 -3 16 105
use FILL  FILL_29
timestamp 1714281807
transform 1 0 2240 0 -1 2970
box -8 -3 16 105
use FILL  FILL_30
timestamp 1714281807
transform 1 0 2232 0 -1 2970
box -8 -3 16 105
use FILL  FILL_31
timestamp 1714281807
transform 1 0 2224 0 -1 2970
box -8 -3 16 105
use FILL  FILL_32
timestamp 1714281807
transform 1 0 2120 0 -1 2970
box -8 -3 16 105
use FILL  FILL_33
timestamp 1714281807
transform 1 0 2112 0 -1 2970
box -8 -3 16 105
use FILL  FILL_34
timestamp 1714281807
transform 1 0 2080 0 -1 2970
box -8 -3 16 105
use FILL  FILL_35
timestamp 1714281807
transform 1 0 2072 0 -1 2970
box -8 -3 16 105
use FILL  FILL_36
timestamp 1714281807
transform 1 0 1872 0 -1 2970
box -8 -3 16 105
use FILL  FILL_37
timestamp 1714281807
transform 1 0 1864 0 -1 2970
box -8 -3 16 105
use FILL  FILL_38
timestamp 1714281807
transform 1 0 1832 0 -1 2970
box -8 -3 16 105
use FILL  FILL_39
timestamp 1714281807
transform 1 0 1824 0 -1 2970
box -8 -3 16 105
use FILL  FILL_40
timestamp 1714281807
transform 1 0 1816 0 -1 2970
box -8 -3 16 105
use FILL  FILL_41
timestamp 1714281807
transform 1 0 1808 0 -1 2970
box -8 -3 16 105
use FILL  FILL_42
timestamp 1714281807
transform 1 0 1776 0 -1 2970
box -8 -3 16 105
use FILL  FILL_43
timestamp 1714281807
transform 1 0 1768 0 -1 2970
box -8 -3 16 105
use FILL  FILL_44
timestamp 1714281807
transform 1 0 1760 0 -1 2970
box -8 -3 16 105
use FILL  FILL_45
timestamp 1714281807
transform 1 0 1560 0 -1 2970
box -8 -3 16 105
use FILL  FILL_46
timestamp 1714281807
transform 1 0 1552 0 -1 2970
box -8 -3 16 105
use FILL  FILL_47
timestamp 1714281807
transform 1 0 1544 0 -1 2970
box -8 -3 16 105
use FILL  FILL_48
timestamp 1714281807
transform 1 0 1512 0 -1 2970
box -8 -3 16 105
use FILL  FILL_49
timestamp 1714281807
transform 1 0 1504 0 -1 2970
box -8 -3 16 105
use FILL  FILL_50
timestamp 1714281807
transform 1 0 1496 0 -1 2970
box -8 -3 16 105
use FILL  FILL_51
timestamp 1714281807
transform 1 0 1472 0 -1 2970
box -8 -3 16 105
use FILL  FILL_52
timestamp 1714281807
transform 1 0 1368 0 -1 2970
box -8 -3 16 105
use FILL  FILL_53
timestamp 1714281807
transform 1 0 1264 0 -1 2970
box -8 -3 16 105
use FILL  FILL_54
timestamp 1714281807
transform 1 0 1256 0 -1 2970
box -8 -3 16 105
use FILL  FILL_55
timestamp 1714281807
transform 1 0 1248 0 -1 2970
box -8 -3 16 105
use FILL  FILL_56
timestamp 1714281807
transform 1 0 1240 0 -1 2970
box -8 -3 16 105
use FILL  FILL_57
timestamp 1714281807
transform 1 0 1232 0 -1 2970
box -8 -3 16 105
use FILL  FILL_58
timestamp 1714281807
transform 1 0 1224 0 -1 2970
box -8 -3 16 105
use FILL  FILL_59
timestamp 1714281807
transform 1 0 1216 0 -1 2970
box -8 -3 16 105
use FILL  FILL_60
timestamp 1714281807
transform 1 0 1208 0 -1 2970
box -8 -3 16 105
use FILL  FILL_61
timestamp 1714281807
transform 1 0 1200 0 -1 2970
box -8 -3 16 105
use FILL  FILL_62
timestamp 1714281807
transform 1 0 1192 0 -1 2970
box -8 -3 16 105
use FILL  FILL_63
timestamp 1714281807
transform 1 0 1184 0 -1 2970
box -8 -3 16 105
use FILL  FILL_64
timestamp 1714281807
transform 1 0 1176 0 -1 2970
box -8 -3 16 105
use FILL  FILL_65
timestamp 1714281807
transform 1 0 1168 0 -1 2970
box -8 -3 16 105
use FILL  FILL_66
timestamp 1714281807
transform 1 0 952 0 -1 2970
box -8 -3 16 105
use FILL  FILL_67
timestamp 1714281807
transform 1 0 888 0 -1 2970
box -8 -3 16 105
use FILL  FILL_68
timestamp 1714281807
transform 1 0 848 0 -1 2970
box -8 -3 16 105
use FILL  FILL_69
timestamp 1714281807
transform 1 0 840 0 -1 2970
box -8 -3 16 105
use FILL  FILL_70
timestamp 1714281807
transform 1 0 736 0 -1 2970
box -8 -3 16 105
use FILL  FILL_71
timestamp 1714281807
transform 1 0 728 0 -1 2970
box -8 -3 16 105
use FILL  FILL_72
timestamp 1714281807
transform 1 0 688 0 -1 2970
box -8 -3 16 105
use FILL  FILL_73
timestamp 1714281807
transform 1 0 680 0 -1 2970
box -8 -3 16 105
use FILL  FILL_74
timestamp 1714281807
transform 1 0 640 0 -1 2970
box -8 -3 16 105
use FILL  FILL_75
timestamp 1714281807
transform 1 0 536 0 -1 2970
box -8 -3 16 105
use FILL  FILL_76
timestamp 1714281807
transform 1 0 528 0 -1 2970
box -8 -3 16 105
use FILL  FILL_77
timestamp 1714281807
transform 1 0 488 0 -1 2970
box -8 -3 16 105
use FILL  FILL_78
timestamp 1714281807
transform 1 0 480 0 -1 2970
box -8 -3 16 105
use FILL  FILL_79
timestamp 1714281807
transform 1 0 472 0 -1 2970
box -8 -3 16 105
use FILL  FILL_80
timestamp 1714281807
transform 1 0 432 0 -1 2970
box -8 -3 16 105
use FILL  FILL_81
timestamp 1714281807
transform 1 0 424 0 -1 2970
box -8 -3 16 105
use FILL  FILL_82
timestamp 1714281807
transform 1 0 416 0 -1 2970
box -8 -3 16 105
use FILL  FILL_83
timestamp 1714281807
transform 1 0 312 0 -1 2970
box -8 -3 16 105
use FILL  FILL_84
timestamp 1714281807
transform 1 0 304 0 -1 2970
box -8 -3 16 105
use FILL  FILL_85
timestamp 1714281807
transform 1 0 296 0 -1 2970
box -8 -3 16 105
use FILL  FILL_86
timestamp 1714281807
transform 1 0 256 0 -1 2970
box -8 -3 16 105
use FILL  FILL_87
timestamp 1714281807
transform 1 0 232 0 -1 2970
box -8 -3 16 105
use FILL  FILL_88
timestamp 1714281807
transform 1 0 224 0 -1 2970
box -8 -3 16 105
use FILL  FILL_89
timestamp 1714281807
transform 1 0 216 0 -1 2970
box -8 -3 16 105
use FILL  FILL_90
timestamp 1714281807
transform 1 0 112 0 -1 2970
box -8 -3 16 105
use FILL  FILL_91
timestamp 1714281807
transform 1 0 104 0 -1 2970
box -8 -3 16 105
use FILL  FILL_92
timestamp 1714281807
transform 1 0 96 0 -1 2970
box -8 -3 16 105
use FILL  FILL_93
timestamp 1714281807
transform 1 0 88 0 -1 2970
box -8 -3 16 105
use FILL  FILL_94
timestamp 1714281807
transform 1 0 80 0 -1 2970
box -8 -3 16 105
use FILL  FILL_95
timestamp 1714281807
transform 1 0 72 0 -1 2970
box -8 -3 16 105
use FILL  FILL_96
timestamp 1714281807
transform 1 0 3000 0 1 2770
box -8 -3 16 105
use FILL  FILL_97
timestamp 1714281807
transform 1 0 2992 0 1 2770
box -8 -3 16 105
use FILL  FILL_98
timestamp 1714281807
transform 1 0 2984 0 1 2770
box -8 -3 16 105
use FILL  FILL_99
timestamp 1714281807
transform 1 0 2976 0 1 2770
box -8 -3 16 105
use FILL  FILL_100
timestamp 1714281807
transform 1 0 2968 0 1 2770
box -8 -3 16 105
use FILL  FILL_101
timestamp 1714281807
transform 1 0 2960 0 1 2770
box -8 -3 16 105
use FILL  FILL_102
timestamp 1714281807
transform 1 0 2952 0 1 2770
box -8 -3 16 105
use FILL  FILL_103
timestamp 1714281807
transform 1 0 2944 0 1 2770
box -8 -3 16 105
use FILL  FILL_104
timestamp 1714281807
transform 1 0 2936 0 1 2770
box -8 -3 16 105
use FILL  FILL_105
timestamp 1714281807
transform 1 0 2928 0 1 2770
box -8 -3 16 105
use FILL  FILL_106
timestamp 1714281807
transform 1 0 2920 0 1 2770
box -8 -3 16 105
use FILL  FILL_107
timestamp 1714281807
transform 1 0 2912 0 1 2770
box -8 -3 16 105
use FILL  FILL_108
timestamp 1714281807
transform 1 0 2904 0 1 2770
box -8 -3 16 105
use FILL  FILL_109
timestamp 1714281807
transform 1 0 2896 0 1 2770
box -8 -3 16 105
use FILL  FILL_110
timestamp 1714281807
transform 1 0 2864 0 1 2770
box -8 -3 16 105
use FILL  FILL_111
timestamp 1714281807
transform 1 0 2856 0 1 2770
box -8 -3 16 105
use FILL  FILL_112
timestamp 1714281807
transform 1 0 2848 0 1 2770
box -8 -3 16 105
use FILL  FILL_113
timestamp 1714281807
transform 1 0 2744 0 1 2770
box -8 -3 16 105
use FILL  FILL_114
timestamp 1714281807
transform 1 0 2736 0 1 2770
box -8 -3 16 105
use FILL  FILL_115
timestamp 1714281807
transform 1 0 2712 0 1 2770
box -8 -3 16 105
use FILL  FILL_116
timestamp 1714281807
transform 1 0 2680 0 1 2770
box -8 -3 16 105
use FILL  FILL_117
timestamp 1714281807
transform 1 0 2672 0 1 2770
box -8 -3 16 105
use FILL  FILL_118
timestamp 1714281807
transform 1 0 2664 0 1 2770
box -8 -3 16 105
use FILL  FILL_119
timestamp 1714281807
transform 1 0 2656 0 1 2770
box -8 -3 16 105
use FILL  FILL_120
timestamp 1714281807
transform 1 0 2648 0 1 2770
box -8 -3 16 105
use FILL  FILL_121
timestamp 1714281807
transform 1 0 2640 0 1 2770
box -8 -3 16 105
use FILL  FILL_122
timestamp 1714281807
transform 1 0 2608 0 1 2770
box -8 -3 16 105
use FILL  FILL_123
timestamp 1714281807
transform 1 0 2600 0 1 2770
box -8 -3 16 105
use FILL  FILL_124
timestamp 1714281807
transform 1 0 2576 0 1 2770
box -8 -3 16 105
use FILL  FILL_125
timestamp 1714281807
transform 1 0 2472 0 1 2770
box -8 -3 16 105
use FILL  FILL_126
timestamp 1714281807
transform 1 0 2352 0 1 2770
box -8 -3 16 105
use FILL  FILL_127
timestamp 1714281807
transform 1 0 2344 0 1 2770
box -8 -3 16 105
use FILL  FILL_128
timestamp 1714281807
transform 1 0 2224 0 1 2770
box -8 -3 16 105
use FILL  FILL_129
timestamp 1714281807
transform 1 0 2216 0 1 2770
box -8 -3 16 105
use FILL  FILL_130
timestamp 1714281807
transform 1 0 2096 0 1 2770
box -8 -3 16 105
use FILL  FILL_131
timestamp 1714281807
transform 1 0 2088 0 1 2770
box -8 -3 16 105
use FILL  FILL_132
timestamp 1714281807
transform 1 0 2080 0 1 2770
box -8 -3 16 105
use FILL  FILL_133
timestamp 1714281807
transform 1 0 2072 0 1 2770
box -8 -3 16 105
use FILL  FILL_134
timestamp 1714281807
transform 1 0 2040 0 1 2770
box -8 -3 16 105
use FILL  FILL_135
timestamp 1714281807
transform 1 0 2032 0 1 2770
box -8 -3 16 105
use FILL  FILL_136
timestamp 1714281807
transform 1 0 1592 0 1 2770
box -8 -3 16 105
use FILL  FILL_137
timestamp 1714281807
transform 1 0 1584 0 1 2770
box -8 -3 16 105
use FILL  FILL_138
timestamp 1714281807
transform 1 0 1552 0 1 2770
box -8 -3 16 105
use FILL  FILL_139
timestamp 1714281807
transform 1 0 1488 0 1 2770
box -8 -3 16 105
use FILL  FILL_140
timestamp 1714281807
transform 1 0 1480 0 1 2770
box -8 -3 16 105
use FILL  FILL_141
timestamp 1714281807
transform 1 0 1472 0 1 2770
box -8 -3 16 105
use FILL  FILL_142
timestamp 1714281807
transform 1 0 1432 0 1 2770
box -8 -3 16 105
use FILL  FILL_143
timestamp 1714281807
transform 1 0 1424 0 1 2770
box -8 -3 16 105
use FILL  FILL_144
timestamp 1714281807
transform 1 0 1416 0 1 2770
box -8 -3 16 105
use FILL  FILL_145
timestamp 1714281807
transform 1 0 1408 0 1 2770
box -8 -3 16 105
use FILL  FILL_146
timestamp 1714281807
transform 1 0 1400 0 1 2770
box -8 -3 16 105
use FILL  FILL_147
timestamp 1714281807
transform 1 0 1392 0 1 2770
box -8 -3 16 105
use FILL  FILL_148
timestamp 1714281807
transform 1 0 1336 0 1 2770
box -8 -3 16 105
use FILL  FILL_149
timestamp 1714281807
transform 1 0 1328 0 1 2770
box -8 -3 16 105
use FILL  FILL_150
timestamp 1714281807
transform 1 0 1320 0 1 2770
box -8 -3 16 105
use FILL  FILL_151
timestamp 1714281807
transform 1 0 1312 0 1 2770
box -8 -3 16 105
use FILL  FILL_152
timestamp 1714281807
transform 1 0 1192 0 1 2770
box -8 -3 16 105
use FILL  FILL_153
timestamp 1714281807
transform 1 0 1184 0 1 2770
box -8 -3 16 105
use FILL  FILL_154
timestamp 1714281807
transform 1 0 1136 0 1 2770
box -8 -3 16 105
use FILL  FILL_155
timestamp 1714281807
transform 1 0 1128 0 1 2770
box -8 -3 16 105
use FILL  FILL_156
timestamp 1714281807
transform 1 0 1120 0 1 2770
box -8 -3 16 105
use FILL  FILL_157
timestamp 1714281807
transform 1 0 1112 0 1 2770
box -8 -3 16 105
use FILL  FILL_158
timestamp 1714281807
transform 1 0 1104 0 1 2770
box -8 -3 16 105
use FILL  FILL_159
timestamp 1714281807
transform 1 0 1056 0 1 2770
box -8 -3 16 105
use FILL  FILL_160
timestamp 1714281807
transform 1 0 1048 0 1 2770
box -8 -3 16 105
use FILL  FILL_161
timestamp 1714281807
transform 1 0 1040 0 1 2770
box -8 -3 16 105
use FILL  FILL_162
timestamp 1714281807
transform 1 0 1032 0 1 2770
box -8 -3 16 105
use FILL  FILL_163
timestamp 1714281807
transform 1 0 1024 0 1 2770
box -8 -3 16 105
use FILL  FILL_164
timestamp 1714281807
transform 1 0 1000 0 1 2770
box -8 -3 16 105
use FILL  FILL_165
timestamp 1714281807
transform 1 0 992 0 1 2770
box -8 -3 16 105
use FILL  FILL_166
timestamp 1714281807
transform 1 0 984 0 1 2770
box -8 -3 16 105
use FILL  FILL_167
timestamp 1714281807
transform 1 0 936 0 1 2770
box -8 -3 16 105
use FILL  FILL_168
timestamp 1714281807
transform 1 0 928 0 1 2770
box -8 -3 16 105
use FILL  FILL_169
timestamp 1714281807
transform 1 0 920 0 1 2770
box -8 -3 16 105
use FILL  FILL_170
timestamp 1714281807
transform 1 0 856 0 1 2770
box -8 -3 16 105
use FILL  FILL_171
timestamp 1714281807
transform 1 0 848 0 1 2770
box -8 -3 16 105
use FILL  FILL_172
timestamp 1714281807
transform 1 0 840 0 1 2770
box -8 -3 16 105
use FILL  FILL_173
timestamp 1714281807
transform 1 0 800 0 1 2770
box -8 -3 16 105
use FILL  FILL_174
timestamp 1714281807
transform 1 0 792 0 1 2770
box -8 -3 16 105
use FILL  FILL_175
timestamp 1714281807
transform 1 0 784 0 1 2770
box -8 -3 16 105
use FILL  FILL_176
timestamp 1714281807
transform 1 0 776 0 1 2770
box -8 -3 16 105
use FILL  FILL_177
timestamp 1714281807
transform 1 0 752 0 1 2770
box -8 -3 16 105
use FILL  FILL_178
timestamp 1714281807
transform 1 0 744 0 1 2770
box -8 -3 16 105
use FILL  FILL_179
timestamp 1714281807
transform 1 0 736 0 1 2770
box -8 -3 16 105
use FILL  FILL_180
timestamp 1714281807
transform 1 0 672 0 1 2770
box -8 -3 16 105
use FILL  FILL_181
timestamp 1714281807
transform 1 0 664 0 1 2770
box -8 -3 16 105
use FILL  FILL_182
timestamp 1714281807
transform 1 0 656 0 1 2770
box -8 -3 16 105
use FILL  FILL_183
timestamp 1714281807
transform 1 0 648 0 1 2770
box -8 -3 16 105
use FILL  FILL_184
timestamp 1714281807
transform 1 0 640 0 1 2770
box -8 -3 16 105
use FILL  FILL_185
timestamp 1714281807
transform 1 0 616 0 1 2770
box -8 -3 16 105
use FILL  FILL_186
timestamp 1714281807
transform 1 0 608 0 1 2770
box -8 -3 16 105
use FILL  FILL_187
timestamp 1714281807
transform 1 0 600 0 1 2770
box -8 -3 16 105
use FILL  FILL_188
timestamp 1714281807
transform 1 0 576 0 1 2770
box -8 -3 16 105
use FILL  FILL_189
timestamp 1714281807
transform 1 0 568 0 1 2770
box -8 -3 16 105
use FILL  FILL_190
timestamp 1714281807
transform 1 0 560 0 1 2770
box -8 -3 16 105
use FILL  FILL_191
timestamp 1714281807
transform 1 0 536 0 1 2770
box -8 -3 16 105
use FILL  FILL_192
timestamp 1714281807
transform 1 0 528 0 1 2770
box -8 -3 16 105
use FILL  FILL_193
timestamp 1714281807
transform 1 0 520 0 1 2770
box -8 -3 16 105
use FILL  FILL_194
timestamp 1714281807
transform 1 0 512 0 1 2770
box -8 -3 16 105
use FILL  FILL_195
timestamp 1714281807
transform 1 0 504 0 1 2770
box -8 -3 16 105
use FILL  FILL_196
timestamp 1714281807
transform 1 0 496 0 1 2770
box -8 -3 16 105
use FILL  FILL_197
timestamp 1714281807
transform 1 0 488 0 1 2770
box -8 -3 16 105
use FILL  FILL_198
timestamp 1714281807
transform 1 0 480 0 1 2770
box -8 -3 16 105
use FILL  FILL_199
timestamp 1714281807
transform 1 0 472 0 1 2770
box -8 -3 16 105
use FILL  FILL_200
timestamp 1714281807
transform 1 0 464 0 1 2770
box -8 -3 16 105
use FILL  FILL_201
timestamp 1714281807
transform 1 0 456 0 1 2770
box -8 -3 16 105
use FILL  FILL_202
timestamp 1714281807
transform 1 0 400 0 1 2770
box -8 -3 16 105
use FILL  FILL_203
timestamp 1714281807
transform 1 0 392 0 1 2770
box -8 -3 16 105
use FILL  FILL_204
timestamp 1714281807
transform 1 0 384 0 1 2770
box -8 -3 16 105
use FILL  FILL_205
timestamp 1714281807
transform 1 0 376 0 1 2770
box -8 -3 16 105
use FILL  FILL_206
timestamp 1714281807
transform 1 0 368 0 1 2770
box -8 -3 16 105
use FILL  FILL_207
timestamp 1714281807
transform 1 0 360 0 1 2770
box -8 -3 16 105
use FILL  FILL_208
timestamp 1714281807
transform 1 0 352 0 1 2770
box -8 -3 16 105
use FILL  FILL_209
timestamp 1714281807
transform 1 0 344 0 1 2770
box -8 -3 16 105
use FILL  FILL_210
timestamp 1714281807
transform 1 0 336 0 1 2770
box -8 -3 16 105
use FILL  FILL_211
timestamp 1714281807
transform 1 0 328 0 1 2770
box -8 -3 16 105
use FILL  FILL_212
timestamp 1714281807
transform 1 0 320 0 1 2770
box -8 -3 16 105
use FILL  FILL_213
timestamp 1714281807
transform 1 0 312 0 1 2770
box -8 -3 16 105
use FILL  FILL_214
timestamp 1714281807
transform 1 0 288 0 1 2770
box -8 -3 16 105
use FILL  FILL_215
timestamp 1714281807
transform 1 0 280 0 1 2770
box -8 -3 16 105
use FILL  FILL_216
timestamp 1714281807
transform 1 0 176 0 1 2770
box -8 -3 16 105
use FILL  FILL_217
timestamp 1714281807
transform 1 0 168 0 1 2770
box -8 -3 16 105
use FILL  FILL_218
timestamp 1714281807
transform 1 0 160 0 1 2770
box -8 -3 16 105
use FILL  FILL_219
timestamp 1714281807
transform 1 0 152 0 1 2770
box -8 -3 16 105
use FILL  FILL_220
timestamp 1714281807
transform 1 0 144 0 1 2770
box -8 -3 16 105
use FILL  FILL_221
timestamp 1714281807
transform 1 0 136 0 1 2770
box -8 -3 16 105
use FILL  FILL_222
timestamp 1714281807
transform 1 0 128 0 1 2770
box -8 -3 16 105
use FILL  FILL_223
timestamp 1714281807
transform 1 0 120 0 1 2770
box -8 -3 16 105
use FILL  FILL_224
timestamp 1714281807
transform 1 0 112 0 1 2770
box -8 -3 16 105
use FILL  FILL_225
timestamp 1714281807
transform 1 0 104 0 1 2770
box -8 -3 16 105
use FILL  FILL_226
timestamp 1714281807
transform 1 0 96 0 1 2770
box -8 -3 16 105
use FILL  FILL_227
timestamp 1714281807
transform 1 0 88 0 1 2770
box -8 -3 16 105
use FILL  FILL_228
timestamp 1714281807
transform 1 0 80 0 1 2770
box -8 -3 16 105
use FILL  FILL_229
timestamp 1714281807
transform 1 0 72 0 1 2770
box -8 -3 16 105
use FILL  FILL_230
timestamp 1714281807
transform 1 0 3000 0 -1 2770
box -8 -3 16 105
use FILL  FILL_231
timestamp 1714281807
transform 1 0 2992 0 -1 2770
box -8 -3 16 105
use FILL  FILL_232
timestamp 1714281807
transform 1 0 2984 0 -1 2770
box -8 -3 16 105
use FILL  FILL_233
timestamp 1714281807
transform 1 0 2976 0 -1 2770
box -8 -3 16 105
use FILL  FILL_234
timestamp 1714281807
transform 1 0 2872 0 -1 2770
box -8 -3 16 105
use FILL  FILL_235
timestamp 1714281807
transform 1 0 2848 0 -1 2770
box -8 -3 16 105
use FILL  FILL_236
timestamp 1714281807
transform 1 0 2840 0 -1 2770
box -8 -3 16 105
use FILL  FILL_237
timestamp 1714281807
transform 1 0 2832 0 -1 2770
box -8 -3 16 105
use FILL  FILL_238
timestamp 1714281807
transform 1 0 2792 0 -1 2770
box -8 -3 16 105
use FILL  FILL_239
timestamp 1714281807
transform 1 0 2784 0 -1 2770
box -8 -3 16 105
use FILL  FILL_240
timestamp 1714281807
transform 1 0 2776 0 -1 2770
box -8 -3 16 105
use FILL  FILL_241
timestamp 1714281807
transform 1 0 2768 0 -1 2770
box -8 -3 16 105
use FILL  FILL_242
timestamp 1714281807
transform 1 0 2760 0 -1 2770
box -8 -3 16 105
use FILL  FILL_243
timestamp 1714281807
transform 1 0 2752 0 -1 2770
box -8 -3 16 105
use FILL  FILL_244
timestamp 1714281807
transform 1 0 2712 0 -1 2770
box -8 -3 16 105
use FILL  FILL_245
timestamp 1714281807
transform 1 0 2704 0 -1 2770
box -8 -3 16 105
use FILL  FILL_246
timestamp 1714281807
transform 1 0 2696 0 -1 2770
box -8 -3 16 105
use FILL  FILL_247
timestamp 1714281807
transform 1 0 2688 0 -1 2770
box -8 -3 16 105
use FILL  FILL_248
timestamp 1714281807
transform 1 0 2624 0 -1 2770
box -8 -3 16 105
use FILL  FILL_249
timestamp 1714281807
transform 1 0 2560 0 -1 2770
box -8 -3 16 105
use FILL  FILL_250
timestamp 1714281807
transform 1 0 2552 0 -1 2770
box -8 -3 16 105
use FILL  FILL_251
timestamp 1714281807
transform 1 0 2544 0 -1 2770
box -8 -3 16 105
use FILL  FILL_252
timestamp 1714281807
transform 1 0 2536 0 -1 2770
box -8 -3 16 105
use FILL  FILL_253
timestamp 1714281807
transform 1 0 2496 0 -1 2770
box -8 -3 16 105
use FILL  FILL_254
timestamp 1714281807
transform 1 0 2488 0 -1 2770
box -8 -3 16 105
use FILL  FILL_255
timestamp 1714281807
transform 1 0 2480 0 -1 2770
box -8 -3 16 105
use FILL  FILL_256
timestamp 1714281807
transform 1 0 2472 0 -1 2770
box -8 -3 16 105
use FILL  FILL_257
timestamp 1714281807
transform 1 0 2464 0 -1 2770
box -8 -3 16 105
use FILL  FILL_258
timestamp 1714281807
transform 1 0 2456 0 -1 2770
box -8 -3 16 105
use FILL  FILL_259
timestamp 1714281807
transform 1 0 2448 0 -1 2770
box -8 -3 16 105
use FILL  FILL_260
timestamp 1714281807
transform 1 0 2408 0 -1 2770
box -8 -3 16 105
use FILL  FILL_261
timestamp 1714281807
transform 1 0 2400 0 -1 2770
box -8 -3 16 105
use FILL  FILL_262
timestamp 1714281807
transform 1 0 2336 0 -1 2770
box -8 -3 16 105
use FILL  FILL_263
timestamp 1714281807
transform 1 0 2328 0 -1 2770
box -8 -3 16 105
use FILL  FILL_264
timestamp 1714281807
transform 1 0 2320 0 -1 2770
box -8 -3 16 105
use FILL  FILL_265
timestamp 1714281807
transform 1 0 2280 0 -1 2770
box -8 -3 16 105
use FILL  FILL_266
timestamp 1714281807
transform 1 0 2272 0 -1 2770
box -8 -3 16 105
use FILL  FILL_267
timestamp 1714281807
transform 1 0 2208 0 -1 2770
box -8 -3 16 105
use FILL  FILL_268
timestamp 1714281807
transform 1 0 2168 0 -1 2770
box -8 -3 16 105
use FILL  FILL_269
timestamp 1714281807
transform 1 0 2160 0 -1 2770
box -8 -3 16 105
use FILL  FILL_270
timestamp 1714281807
transform 1 0 2152 0 -1 2770
box -8 -3 16 105
use FILL  FILL_271
timestamp 1714281807
transform 1 0 2088 0 -1 2770
box -8 -3 16 105
use FILL  FILL_272
timestamp 1714281807
transform 1 0 2048 0 -1 2770
box -8 -3 16 105
use FILL  FILL_273
timestamp 1714281807
transform 1 0 2040 0 -1 2770
box -8 -3 16 105
use FILL  FILL_274
timestamp 1714281807
transform 1 0 2032 0 -1 2770
box -8 -3 16 105
use FILL  FILL_275
timestamp 1714281807
transform 1 0 2024 0 -1 2770
box -8 -3 16 105
use FILL  FILL_276
timestamp 1714281807
transform 1 0 2016 0 -1 2770
box -8 -3 16 105
use FILL  FILL_277
timestamp 1714281807
transform 1 0 2008 0 -1 2770
box -8 -3 16 105
use FILL  FILL_278
timestamp 1714281807
transform 1 0 2000 0 -1 2770
box -8 -3 16 105
use FILL  FILL_279
timestamp 1714281807
transform 1 0 1992 0 -1 2770
box -8 -3 16 105
use FILL  FILL_280
timestamp 1714281807
transform 1 0 1952 0 -1 2770
box -8 -3 16 105
use FILL  FILL_281
timestamp 1714281807
transform 1 0 1944 0 -1 2770
box -8 -3 16 105
use FILL  FILL_282
timestamp 1714281807
transform 1 0 1936 0 -1 2770
box -8 -3 16 105
use FILL  FILL_283
timestamp 1714281807
transform 1 0 1928 0 -1 2770
box -8 -3 16 105
use FILL  FILL_284
timestamp 1714281807
transform 1 0 1920 0 -1 2770
box -8 -3 16 105
use FILL  FILL_285
timestamp 1714281807
transform 1 0 1912 0 -1 2770
box -8 -3 16 105
use FILL  FILL_286
timestamp 1714281807
transform 1 0 1904 0 -1 2770
box -8 -3 16 105
use FILL  FILL_287
timestamp 1714281807
transform 1 0 1864 0 -1 2770
box -8 -3 16 105
use FILL  FILL_288
timestamp 1714281807
transform 1 0 1856 0 -1 2770
box -8 -3 16 105
use FILL  FILL_289
timestamp 1714281807
transform 1 0 1792 0 -1 2770
box -8 -3 16 105
use FILL  FILL_290
timestamp 1714281807
transform 1 0 1752 0 -1 2770
box -8 -3 16 105
use FILL  FILL_291
timestamp 1714281807
transform 1 0 1744 0 -1 2770
box -8 -3 16 105
use FILL  FILL_292
timestamp 1714281807
transform 1 0 1640 0 -1 2770
box -8 -3 16 105
use FILL  FILL_293
timestamp 1714281807
transform 1 0 1608 0 -1 2770
box -8 -3 16 105
use FILL  FILL_294
timestamp 1714281807
transform 1 0 1600 0 -1 2770
box -8 -3 16 105
use FILL  FILL_295
timestamp 1714281807
transform 1 0 1560 0 -1 2770
box -8 -3 16 105
use FILL  FILL_296
timestamp 1714281807
transform 1 0 1496 0 -1 2770
box -8 -3 16 105
use FILL  FILL_297
timestamp 1714281807
transform 1 0 1448 0 -1 2770
box -8 -3 16 105
use FILL  FILL_298
timestamp 1714281807
transform 1 0 1440 0 -1 2770
box -8 -3 16 105
use FILL  FILL_299
timestamp 1714281807
transform 1 0 1432 0 -1 2770
box -8 -3 16 105
use FILL  FILL_300
timestamp 1714281807
transform 1 0 1424 0 -1 2770
box -8 -3 16 105
use FILL  FILL_301
timestamp 1714281807
transform 1 0 1376 0 -1 2770
box -8 -3 16 105
use FILL  FILL_302
timestamp 1714281807
transform 1 0 1368 0 -1 2770
box -8 -3 16 105
use FILL  FILL_303
timestamp 1714281807
transform 1 0 984 0 -1 2770
box -8 -3 16 105
use FILL  FILL_304
timestamp 1714281807
transform 1 0 936 0 -1 2770
box -8 -3 16 105
use FILL  FILL_305
timestamp 1714281807
transform 1 0 640 0 -1 2770
box -8 -3 16 105
use FILL  FILL_306
timestamp 1714281807
transform 1 0 600 0 -1 2770
box -8 -3 16 105
use FILL  FILL_307
timestamp 1714281807
transform 1 0 576 0 -1 2770
box -8 -3 16 105
use FILL  FILL_308
timestamp 1714281807
transform 1 0 568 0 -1 2770
box -8 -3 16 105
use FILL  FILL_309
timestamp 1714281807
transform 1 0 424 0 -1 2770
box -8 -3 16 105
use FILL  FILL_310
timestamp 1714281807
transform 1 0 416 0 -1 2770
box -8 -3 16 105
use FILL  FILL_311
timestamp 1714281807
transform 1 0 408 0 -1 2770
box -8 -3 16 105
use FILL  FILL_312
timestamp 1714281807
transform 1 0 344 0 -1 2770
box -8 -3 16 105
use FILL  FILL_313
timestamp 1714281807
transform 1 0 240 0 -1 2770
box -8 -3 16 105
use FILL  FILL_314
timestamp 1714281807
transform 1 0 192 0 -1 2770
box -8 -3 16 105
use FILL  FILL_315
timestamp 1714281807
transform 1 0 184 0 -1 2770
box -8 -3 16 105
use FILL  FILL_316
timestamp 1714281807
transform 1 0 176 0 -1 2770
box -8 -3 16 105
use FILL  FILL_317
timestamp 1714281807
transform 1 0 168 0 -1 2770
box -8 -3 16 105
use FILL  FILL_318
timestamp 1714281807
transform 1 0 160 0 -1 2770
box -8 -3 16 105
use FILL  FILL_319
timestamp 1714281807
transform 1 0 152 0 -1 2770
box -8 -3 16 105
use FILL  FILL_320
timestamp 1714281807
transform 1 0 144 0 -1 2770
box -8 -3 16 105
use FILL  FILL_321
timestamp 1714281807
transform 1 0 136 0 -1 2770
box -8 -3 16 105
use FILL  FILL_322
timestamp 1714281807
transform 1 0 128 0 -1 2770
box -8 -3 16 105
use FILL  FILL_323
timestamp 1714281807
transform 1 0 120 0 -1 2770
box -8 -3 16 105
use FILL  FILL_324
timestamp 1714281807
transform 1 0 112 0 -1 2770
box -8 -3 16 105
use FILL  FILL_325
timestamp 1714281807
transform 1 0 104 0 -1 2770
box -8 -3 16 105
use FILL  FILL_326
timestamp 1714281807
transform 1 0 96 0 -1 2770
box -8 -3 16 105
use FILL  FILL_327
timestamp 1714281807
transform 1 0 88 0 -1 2770
box -8 -3 16 105
use FILL  FILL_328
timestamp 1714281807
transform 1 0 80 0 -1 2770
box -8 -3 16 105
use FILL  FILL_329
timestamp 1714281807
transform 1 0 72 0 -1 2770
box -8 -3 16 105
use FILL  FILL_330
timestamp 1714281807
transform 1 0 3000 0 1 2570
box -8 -3 16 105
use FILL  FILL_331
timestamp 1714281807
transform 1 0 2992 0 1 2570
box -8 -3 16 105
use FILL  FILL_332
timestamp 1714281807
transform 1 0 2984 0 1 2570
box -8 -3 16 105
use FILL  FILL_333
timestamp 1714281807
transform 1 0 2976 0 1 2570
box -8 -3 16 105
use FILL  FILL_334
timestamp 1714281807
transform 1 0 2968 0 1 2570
box -8 -3 16 105
use FILL  FILL_335
timestamp 1714281807
transform 1 0 2960 0 1 2570
box -8 -3 16 105
use FILL  FILL_336
timestamp 1714281807
transform 1 0 2952 0 1 2570
box -8 -3 16 105
use FILL  FILL_337
timestamp 1714281807
transform 1 0 2944 0 1 2570
box -8 -3 16 105
use FILL  FILL_338
timestamp 1714281807
transform 1 0 2936 0 1 2570
box -8 -3 16 105
use FILL  FILL_339
timestamp 1714281807
transform 1 0 2928 0 1 2570
box -8 -3 16 105
use FILL  FILL_340
timestamp 1714281807
transform 1 0 2920 0 1 2570
box -8 -3 16 105
use FILL  FILL_341
timestamp 1714281807
transform 1 0 2912 0 1 2570
box -8 -3 16 105
use FILL  FILL_342
timestamp 1714281807
transform 1 0 2904 0 1 2570
box -8 -3 16 105
use FILL  FILL_343
timestamp 1714281807
transform 1 0 2840 0 1 2570
box -8 -3 16 105
use FILL  FILL_344
timestamp 1714281807
transform 1 0 2832 0 1 2570
box -8 -3 16 105
use FILL  FILL_345
timestamp 1714281807
transform 1 0 2824 0 1 2570
box -8 -3 16 105
use FILL  FILL_346
timestamp 1714281807
transform 1 0 2776 0 1 2570
box -8 -3 16 105
use FILL  FILL_347
timestamp 1714281807
transform 1 0 2768 0 1 2570
box -8 -3 16 105
use FILL  FILL_348
timestamp 1714281807
transform 1 0 2760 0 1 2570
box -8 -3 16 105
use FILL  FILL_349
timestamp 1714281807
transform 1 0 2752 0 1 2570
box -8 -3 16 105
use FILL  FILL_350
timestamp 1714281807
transform 1 0 2744 0 1 2570
box -8 -3 16 105
use FILL  FILL_351
timestamp 1714281807
transform 1 0 2736 0 1 2570
box -8 -3 16 105
use FILL  FILL_352
timestamp 1714281807
transform 1 0 2688 0 1 2570
box -8 -3 16 105
use FILL  FILL_353
timestamp 1714281807
transform 1 0 2680 0 1 2570
box -8 -3 16 105
use FILL  FILL_354
timestamp 1714281807
transform 1 0 2672 0 1 2570
box -8 -3 16 105
use FILL  FILL_355
timestamp 1714281807
transform 1 0 2664 0 1 2570
box -8 -3 16 105
use FILL  FILL_356
timestamp 1714281807
transform 1 0 2656 0 1 2570
box -8 -3 16 105
use FILL  FILL_357
timestamp 1714281807
transform 1 0 2616 0 1 2570
box -8 -3 16 105
use FILL  FILL_358
timestamp 1714281807
transform 1 0 2608 0 1 2570
box -8 -3 16 105
use FILL  FILL_359
timestamp 1714281807
transform 1 0 2600 0 1 2570
box -8 -3 16 105
use FILL  FILL_360
timestamp 1714281807
transform 1 0 2560 0 1 2570
box -8 -3 16 105
use FILL  FILL_361
timestamp 1714281807
transform 1 0 2552 0 1 2570
box -8 -3 16 105
use FILL  FILL_362
timestamp 1714281807
transform 1 0 2544 0 1 2570
box -8 -3 16 105
use FILL  FILL_363
timestamp 1714281807
transform 1 0 2496 0 1 2570
box -8 -3 16 105
use FILL  FILL_364
timestamp 1714281807
transform 1 0 2488 0 1 2570
box -8 -3 16 105
use FILL  FILL_365
timestamp 1714281807
transform 1 0 2480 0 1 2570
box -8 -3 16 105
use FILL  FILL_366
timestamp 1714281807
transform 1 0 2472 0 1 2570
box -8 -3 16 105
use FILL  FILL_367
timestamp 1714281807
transform 1 0 2464 0 1 2570
box -8 -3 16 105
use FILL  FILL_368
timestamp 1714281807
transform 1 0 2456 0 1 2570
box -8 -3 16 105
use FILL  FILL_369
timestamp 1714281807
transform 1 0 2424 0 1 2570
box -8 -3 16 105
use FILL  FILL_370
timestamp 1714281807
transform 1 0 2416 0 1 2570
box -8 -3 16 105
use FILL  FILL_371
timestamp 1714281807
transform 1 0 2408 0 1 2570
box -8 -3 16 105
use FILL  FILL_372
timestamp 1714281807
transform 1 0 2360 0 1 2570
box -8 -3 16 105
use FILL  FILL_373
timestamp 1714281807
transform 1 0 2352 0 1 2570
box -8 -3 16 105
use FILL  FILL_374
timestamp 1714281807
transform 1 0 2344 0 1 2570
box -8 -3 16 105
use FILL  FILL_375
timestamp 1714281807
transform 1 0 2336 0 1 2570
box -8 -3 16 105
use FILL  FILL_376
timestamp 1714281807
transform 1 0 2328 0 1 2570
box -8 -3 16 105
use FILL  FILL_377
timestamp 1714281807
transform 1 0 2320 0 1 2570
box -8 -3 16 105
use FILL  FILL_378
timestamp 1714281807
transform 1 0 2272 0 1 2570
box -8 -3 16 105
use FILL  FILL_379
timestamp 1714281807
transform 1 0 2264 0 1 2570
box -8 -3 16 105
use FILL  FILL_380
timestamp 1714281807
transform 1 0 2256 0 1 2570
box -8 -3 16 105
use FILL  FILL_381
timestamp 1714281807
transform 1 0 2248 0 1 2570
box -8 -3 16 105
use FILL  FILL_382
timestamp 1714281807
transform 1 0 2208 0 1 2570
box -8 -3 16 105
use FILL  FILL_383
timestamp 1714281807
transform 1 0 2200 0 1 2570
box -8 -3 16 105
use FILL  FILL_384
timestamp 1714281807
transform 1 0 2168 0 1 2570
box -8 -3 16 105
use FILL  FILL_385
timestamp 1714281807
transform 1 0 2160 0 1 2570
box -8 -3 16 105
use FILL  FILL_386
timestamp 1714281807
transform 1 0 2152 0 1 2570
box -8 -3 16 105
use FILL  FILL_387
timestamp 1714281807
transform 1 0 2144 0 1 2570
box -8 -3 16 105
use FILL  FILL_388
timestamp 1714281807
transform 1 0 2136 0 1 2570
box -8 -3 16 105
use FILL  FILL_389
timestamp 1714281807
transform 1 0 2088 0 1 2570
box -8 -3 16 105
use FILL  FILL_390
timestamp 1714281807
transform 1 0 2080 0 1 2570
box -8 -3 16 105
use FILL  FILL_391
timestamp 1714281807
transform 1 0 2072 0 1 2570
box -8 -3 16 105
use FILL  FILL_392
timestamp 1714281807
transform 1 0 2064 0 1 2570
box -8 -3 16 105
use FILL  FILL_393
timestamp 1714281807
transform 1 0 2056 0 1 2570
box -8 -3 16 105
use FILL  FILL_394
timestamp 1714281807
transform 1 0 1960 0 1 2570
box -8 -3 16 105
use FILL  FILL_395
timestamp 1714281807
transform 1 0 1952 0 1 2570
box -8 -3 16 105
use FILL  FILL_396
timestamp 1714281807
transform 1 0 1848 0 1 2570
box -8 -3 16 105
use FILL  FILL_397
timestamp 1714281807
transform 1 0 1840 0 1 2570
box -8 -3 16 105
use FILL  FILL_398
timestamp 1714281807
transform 1 0 1832 0 1 2570
box -8 -3 16 105
use FILL  FILL_399
timestamp 1714281807
transform 1 0 1784 0 1 2570
box -8 -3 16 105
use FILL  FILL_400
timestamp 1714281807
transform 1 0 1776 0 1 2570
box -8 -3 16 105
use FILL  FILL_401
timestamp 1714281807
transform 1 0 1768 0 1 2570
box -8 -3 16 105
use FILL  FILL_402
timestamp 1714281807
transform 1 0 1760 0 1 2570
box -8 -3 16 105
use FILL  FILL_403
timestamp 1714281807
transform 1 0 1752 0 1 2570
box -8 -3 16 105
use FILL  FILL_404
timestamp 1714281807
transform 1 0 1704 0 1 2570
box -8 -3 16 105
use FILL  FILL_405
timestamp 1714281807
transform 1 0 1696 0 1 2570
box -8 -3 16 105
use FILL  FILL_406
timestamp 1714281807
transform 1 0 1688 0 1 2570
box -8 -3 16 105
use FILL  FILL_407
timestamp 1714281807
transform 1 0 1680 0 1 2570
box -8 -3 16 105
use FILL  FILL_408
timestamp 1714281807
transform 1 0 1672 0 1 2570
box -8 -3 16 105
use FILL  FILL_409
timestamp 1714281807
transform 1 0 1632 0 1 2570
box -8 -3 16 105
use FILL  FILL_410
timestamp 1714281807
transform 1 0 1568 0 1 2570
box -8 -3 16 105
use FILL  FILL_411
timestamp 1714281807
transform 1 0 1464 0 1 2570
box -8 -3 16 105
use FILL  FILL_412
timestamp 1714281807
transform 1 0 1456 0 1 2570
box -8 -3 16 105
use FILL  FILL_413
timestamp 1714281807
transform 1 0 1448 0 1 2570
box -8 -3 16 105
use FILL  FILL_414
timestamp 1714281807
transform 1 0 1400 0 1 2570
box -8 -3 16 105
use FILL  FILL_415
timestamp 1714281807
transform 1 0 1392 0 1 2570
box -8 -3 16 105
use FILL  FILL_416
timestamp 1714281807
transform 1 0 1384 0 1 2570
box -8 -3 16 105
use FILL  FILL_417
timestamp 1714281807
transform 1 0 1344 0 1 2570
box -8 -3 16 105
use FILL  FILL_418
timestamp 1714281807
transform 1 0 1336 0 1 2570
box -8 -3 16 105
use FILL  FILL_419
timestamp 1714281807
transform 1 0 1328 0 1 2570
box -8 -3 16 105
use FILL  FILL_420
timestamp 1714281807
transform 1 0 1288 0 1 2570
box -8 -3 16 105
use FILL  FILL_421
timestamp 1714281807
transform 1 0 1280 0 1 2570
box -8 -3 16 105
use FILL  FILL_422
timestamp 1714281807
transform 1 0 1272 0 1 2570
box -8 -3 16 105
use FILL  FILL_423
timestamp 1714281807
transform 1 0 1264 0 1 2570
box -8 -3 16 105
use FILL  FILL_424
timestamp 1714281807
transform 1 0 1256 0 1 2570
box -8 -3 16 105
use FILL  FILL_425
timestamp 1714281807
transform 1 0 1248 0 1 2570
box -8 -3 16 105
use FILL  FILL_426
timestamp 1714281807
transform 1 0 1216 0 1 2570
box -8 -3 16 105
use FILL  FILL_427
timestamp 1714281807
transform 1 0 1208 0 1 2570
box -8 -3 16 105
use FILL  FILL_428
timestamp 1714281807
transform 1 0 1200 0 1 2570
box -8 -3 16 105
use FILL  FILL_429
timestamp 1714281807
transform 1 0 1192 0 1 2570
box -8 -3 16 105
use FILL  FILL_430
timestamp 1714281807
transform 1 0 1160 0 1 2570
box -8 -3 16 105
use FILL  FILL_431
timestamp 1714281807
transform 1 0 1152 0 1 2570
box -8 -3 16 105
use FILL  FILL_432
timestamp 1714281807
transform 1 0 1144 0 1 2570
box -8 -3 16 105
use FILL  FILL_433
timestamp 1714281807
transform 1 0 1136 0 1 2570
box -8 -3 16 105
use FILL  FILL_434
timestamp 1714281807
transform 1 0 1128 0 1 2570
box -8 -3 16 105
use FILL  FILL_435
timestamp 1714281807
transform 1 0 1120 0 1 2570
box -8 -3 16 105
use FILL  FILL_436
timestamp 1714281807
transform 1 0 1112 0 1 2570
box -8 -3 16 105
use FILL  FILL_437
timestamp 1714281807
transform 1 0 1048 0 1 2570
box -8 -3 16 105
use FILL  FILL_438
timestamp 1714281807
transform 1 0 1040 0 1 2570
box -8 -3 16 105
use FILL  FILL_439
timestamp 1714281807
transform 1 0 1032 0 1 2570
box -8 -3 16 105
use FILL  FILL_440
timestamp 1714281807
transform 1 0 928 0 1 2570
box -8 -3 16 105
use FILL  FILL_441
timestamp 1714281807
transform 1 0 920 0 1 2570
box -8 -3 16 105
use FILL  FILL_442
timestamp 1714281807
transform 1 0 912 0 1 2570
box -8 -3 16 105
use FILL  FILL_443
timestamp 1714281807
transform 1 0 904 0 1 2570
box -8 -3 16 105
use FILL  FILL_444
timestamp 1714281807
transform 1 0 840 0 1 2570
box -8 -3 16 105
use FILL  FILL_445
timestamp 1714281807
transform 1 0 832 0 1 2570
box -8 -3 16 105
use FILL  FILL_446
timestamp 1714281807
transform 1 0 824 0 1 2570
box -8 -3 16 105
use FILL  FILL_447
timestamp 1714281807
transform 1 0 816 0 1 2570
box -8 -3 16 105
use FILL  FILL_448
timestamp 1714281807
transform 1 0 808 0 1 2570
box -8 -3 16 105
use FILL  FILL_449
timestamp 1714281807
transform 1 0 800 0 1 2570
box -8 -3 16 105
use FILL  FILL_450
timestamp 1714281807
transform 1 0 752 0 1 2570
box -8 -3 16 105
use FILL  FILL_451
timestamp 1714281807
transform 1 0 728 0 1 2570
box -8 -3 16 105
use FILL  FILL_452
timestamp 1714281807
transform 1 0 720 0 1 2570
box -8 -3 16 105
use FILL  FILL_453
timestamp 1714281807
transform 1 0 712 0 1 2570
box -8 -3 16 105
use FILL  FILL_454
timestamp 1714281807
transform 1 0 704 0 1 2570
box -8 -3 16 105
use FILL  FILL_455
timestamp 1714281807
transform 1 0 584 0 1 2570
box -8 -3 16 105
use FILL  FILL_456
timestamp 1714281807
transform 1 0 576 0 1 2570
box -8 -3 16 105
use FILL  FILL_457
timestamp 1714281807
transform 1 0 528 0 1 2570
box -8 -3 16 105
use FILL  FILL_458
timestamp 1714281807
transform 1 0 520 0 1 2570
box -8 -3 16 105
use FILL  FILL_459
timestamp 1714281807
transform 1 0 512 0 1 2570
box -8 -3 16 105
use FILL  FILL_460
timestamp 1714281807
transform 1 0 504 0 1 2570
box -8 -3 16 105
use FILL  FILL_461
timestamp 1714281807
transform 1 0 496 0 1 2570
box -8 -3 16 105
use FILL  FILL_462
timestamp 1714281807
transform 1 0 488 0 1 2570
box -8 -3 16 105
use FILL  FILL_463
timestamp 1714281807
transform 1 0 480 0 1 2570
box -8 -3 16 105
use FILL  FILL_464
timestamp 1714281807
transform 1 0 416 0 1 2570
box -8 -3 16 105
use FILL  FILL_465
timestamp 1714281807
transform 1 0 312 0 1 2570
box -8 -3 16 105
use FILL  FILL_466
timestamp 1714281807
transform 1 0 304 0 1 2570
box -8 -3 16 105
use FILL  FILL_467
timestamp 1714281807
transform 1 0 296 0 1 2570
box -8 -3 16 105
use FILL  FILL_468
timestamp 1714281807
transform 1 0 288 0 1 2570
box -8 -3 16 105
use FILL  FILL_469
timestamp 1714281807
transform 1 0 240 0 1 2570
box -8 -3 16 105
use FILL  FILL_470
timestamp 1714281807
transform 1 0 232 0 1 2570
box -8 -3 16 105
use FILL  FILL_471
timestamp 1714281807
transform 1 0 224 0 1 2570
box -8 -3 16 105
use FILL  FILL_472
timestamp 1714281807
transform 1 0 216 0 1 2570
box -8 -3 16 105
use FILL  FILL_473
timestamp 1714281807
transform 1 0 208 0 1 2570
box -8 -3 16 105
use FILL  FILL_474
timestamp 1714281807
transform 1 0 88 0 1 2570
box -8 -3 16 105
use FILL  FILL_475
timestamp 1714281807
transform 1 0 80 0 1 2570
box -8 -3 16 105
use FILL  FILL_476
timestamp 1714281807
transform 1 0 72 0 1 2570
box -8 -3 16 105
use FILL  FILL_477
timestamp 1714281807
transform 1 0 3000 0 -1 2570
box -8 -3 16 105
use FILL  FILL_478
timestamp 1714281807
transform 1 0 2992 0 -1 2570
box -8 -3 16 105
use FILL  FILL_479
timestamp 1714281807
transform 1 0 2984 0 -1 2570
box -8 -3 16 105
use FILL  FILL_480
timestamp 1714281807
transform 1 0 2976 0 -1 2570
box -8 -3 16 105
use FILL  FILL_481
timestamp 1714281807
transform 1 0 2968 0 -1 2570
box -8 -3 16 105
use FILL  FILL_482
timestamp 1714281807
transform 1 0 2864 0 -1 2570
box -8 -3 16 105
use FILL  FILL_483
timestamp 1714281807
transform 1 0 2856 0 -1 2570
box -8 -3 16 105
use FILL  FILL_484
timestamp 1714281807
transform 1 0 2848 0 -1 2570
box -8 -3 16 105
use FILL  FILL_485
timestamp 1714281807
transform 1 0 2840 0 -1 2570
box -8 -3 16 105
use FILL  FILL_486
timestamp 1714281807
transform 1 0 2832 0 -1 2570
box -8 -3 16 105
use FILL  FILL_487
timestamp 1714281807
transform 1 0 2784 0 -1 2570
box -8 -3 16 105
use FILL  FILL_488
timestamp 1714281807
transform 1 0 2776 0 -1 2570
box -8 -3 16 105
use FILL  FILL_489
timestamp 1714281807
transform 1 0 2768 0 -1 2570
box -8 -3 16 105
use FILL  FILL_490
timestamp 1714281807
transform 1 0 2760 0 -1 2570
box -8 -3 16 105
use FILL  FILL_491
timestamp 1714281807
transform 1 0 2560 0 -1 2570
box -8 -3 16 105
use FILL  FILL_492
timestamp 1714281807
transform 1 0 2552 0 -1 2570
box -8 -3 16 105
use FILL  FILL_493
timestamp 1714281807
transform 1 0 2528 0 -1 2570
box -8 -3 16 105
use FILL  FILL_494
timestamp 1714281807
transform 1 0 2424 0 -1 2570
box -8 -3 16 105
use FILL  FILL_495
timestamp 1714281807
transform 1 0 2416 0 -1 2570
box -8 -3 16 105
use FILL  FILL_496
timestamp 1714281807
transform 1 0 2408 0 -1 2570
box -8 -3 16 105
use FILL  FILL_497
timestamp 1714281807
transform 1 0 2288 0 -1 2570
box -8 -3 16 105
use FILL  FILL_498
timestamp 1714281807
transform 1 0 2280 0 -1 2570
box -8 -3 16 105
use FILL  FILL_499
timestamp 1714281807
transform 1 0 1952 0 -1 2570
box -8 -3 16 105
use FILL  FILL_500
timestamp 1714281807
transform 1 0 1944 0 -1 2570
box -8 -3 16 105
use FILL  FILL_501
timestamp 1714281807
transform 1 0 1840 0 -1 2570
box -8 -3 16 105
use FILL  FILL_502
timestamp 1714281807
transform 1 0 1720 0 -1 2570
box -8 -3 16 105
use FILL  FILL_503
timestamp 1714281807
transform 1 0 1712 0 -1 2570
box -8 -3 16 105
use FILL  FILL_504
timestamp 1714281807
transform 1 0 1608 0 -1 2570
box -8 -3 16 105
use FILL  FILL_505
timestamp 1714281807
transform 1 0 1600 0 -1 2570
box -8 -3 16 105
use FILL  FILL_506
timestamp 1714281807
transform 1 0 1592 0 -1 2570
box -8 -3 16 105
use FILL  FILL_507
timestamp 1714281807
transform 1 0 1560 0 -1 2570
box -8 -3 16 105
use FILL  FILL_508
timestamp 1714281807
transform 1 0 1552 0 -1 2570
box -8 -3 16 105
use FILL  FILL_509
timestamp 1714281807
transform 1 0 1544 0 -1 2570
box -8 -3 16 105
use FILL  FILL_510
timestamp 1714281807
transform 1 0 1536 0 -1 2570
box -8 -3 16 105
use FILL  FILL_511
timestamp 1714281807
transform 1 0 1496 0 -1 2570
box -8 -3 16 105
use FILL  FILL_512
timestamp 1714281807
transform 1 0 1488 0 -1 2570
box -8 -3 16 105
use FILL  FILL_513
timestamp 1714281807
transform 1 0 1096 0 -1 2570
box -8 -3 16 105
use FILL  FILL_514
timestamp 1714281807
transform 1 0 1088 0 -1 2570
box -8 -3 16 105
use FILL  FILL_515
timestamp 1714281807
transform 1 0 1056 0 -1 2570
box -8 -3 16 105
use FILL  FILL_516
timestamp 1714281807
transform 1 0 1048 0 -1 2570
box -8 -3 16 105
use FILL  FILL_517
timestamp 1714281807
transform 1 0 1040 0 -1 2570
box -8 -3 16 105
use FILL  FILL_518
timestamp 1714281807
transform 1 0 1032 0 -1 2570
box -8 -3 16 105
use FILL  FILL_519
timestamp 1714281807
transform 1 0 1000 0 -1 2570
box -8 -3 16 105
use FILL  FILL_520
timestamp 1714281807
transform 1 0 992 0 -1 2570
box -8 -3 16 105
use FILL  FILL_521
timestamp 1714281807
transform 1 0 984 0 -1 2570
box -8 -3 16 105
use FILL  FILL_522
timestamp 1714281807
transform 1 0 976 0 -1 2570
box -8 -3 16 105
use FILL  FILL_523
timestamp 1714281807
transform 1 0 944 0 -1 2570
box -8 -3 16 105
use FILL  FILL_524
timestamp 1714281807
transform 1 0 936 0 -1 2570
box -8 -3 16 105
use FILL  FILL_525
timestamp 1714281807
transform 1 0 928 0 -1 2570
box -8 -3 16 105
use FILL  FILL_526
timestamp 1714281807
transform 1 0 808 0 -1 2570
box -8 -3 16 105
use FILL  FILL_527
timestamp 1714281807
transform 1 0 800 0 -1 2570
box -8 -3 16 105
use FILL  FILL_528
timestamp 1714281807
transform 1 0 680 0 -1 2570
box -8 -3 16 105
use FILL  FILL_529
timestamp 1714281807
transform 1 0 672 0 -1 2570
box -8 -3 16 105
use FILL  FILL_530
timestamp 1714281807
transform 1 0 664 0 -1 2570
box -8 -3 16 105
use FILL  FILL_531
timestamp 1714281807
transform 1 0 656 0 -1 2570
box -8 -3 16 105
use FILL  FILL_532
timestamp 1714281807
transform 1 0 648 0 -1 2570
box -8 -3 16 105
use FILL  FILL_533
timestamp 1714281807
transform 1 0 640 0 -1 2570
box -8 -3 16 105
use FILL  FILL_534
timestamp 1714281807
transform 1 0 632 0 -1 2570
box -8 -3 16 105
use FILL  FILL_535
timestamp 1714281807
transform 1 0 584 0 -1 2570
box -8 -3 16 105
use FILL  FILL_536
timestamp 1714281807
transform 1 0 576 0 -1 2570
box -8 -3 16 105
use FILL  FILL_537
timestamp 1714281807
transform 1 0 568 0 -1 2570
box -8 -3 16 105
use FILL  FILL_538
timestamp 1714281807
transform 1 0 560 0 -1 2570
box -8 -3 16 105
use FILL  FILL_539
timestamp 1714281807
transform 1 0 552 0 -1 2570
box -8 -3 16 105
use FILL  FILL_540
timestamp 1714281807
transform 1 0 544 0 -1 2570
box -8 -3 16 105
use FILL  FILL_541
timestamp 1714281807
transform 1 0 496 0 -1 2570
box -8 -3 16 105
use FILL  FILL_542
timestamp 1714281807
transform 1 0 488 0 -1 2570
box -8 -3 16 105
use FILL  FILL_543
timestamp 1714281807
transform 1 0 464 0 -1 2570
box -8 -3 16 105
use FILL  FILL_544
timestamp 1714281807
transform 1 0 456 0 -1 2570
box -8 -3 16 105
use FILL  FILL_545
timestamp 1714281807
transform 1 0 352 0 -1 2570
box -8 -3 16 105
use FILL  FILL_546
timestamp 1714281807
transform 1 0 344 0 -1 2570
box -8 -3 16 105
use FILL  FILL_547
timestamp 1714281807
transform 1 0 336 0 -1 2570
box -8 -3 16 105
use FILL  FILL_548
timestamp 1714281807
transform 1 0 328 0 -1 2570
box -8 -3 16 105
use FILL  FILL_549
timestamp 1714281807
transform 1 0 264 0 -1 2570
box -8 -3 16 105
use FILL  FILL_550
timestamp 1714281807
transform 1 0 256 0 -1 2570
box -8 -3 16 105
use FILL  FILL_551
timestamp 1714281807
transform 1 0 248 0 -1 2570
box -8 -3 16 105
use FILL  FILL_552
timestamp 1714281807
transform 1 0 144 0 -1 2570
box -8 -3 16 105
use FILL  FILL_553
timestamp 1714281807
transform 1 0 136 0 -1 2570
box -8 -3 16 105
use FILL  FILL_554
timestamp 1714281807
transform 1 0 128 0 -1 2570
box -8 -3 16 105
use FILL  FILL_555
timestamp 1714281807
transform 1 0 120 0 -1 2570
box -8 -3 16 105
use FILL  FILL_556
timestamp 1714281807
transform 1 0 112 0 -1 2570
box -8 -3 16 105
use FILL  FILL_557
timestamp 1714281807
transform 1 0 104 0 -1 2570
box -8 -3 16 105
use FILL  FILL_558
timestamp 1714281807
transform 1 0 96 0 -1 2570
box -8 -3 16 105
use FILL  FILL_559
timestamp 1714281807
transform 1 0 88 0 -1 2570
box -8 -3 16 105
use FILL  FILL_560
timestamp 1714281807
transform 1 0 80 0 -1 2570
box -8 -3 16 105
use FILL  FILL_561
timestamp 1714281807
transform 1 0 72 0 -1 2570
box -8 -3 16 105
use FILL  FILL_562
timestamp 1714281807
transform 1 0 3000 0 1 2370
box -8 -3 16 105
use FILL  FILL_563
timestamp 1714281807
transform 1 0 2992 0 1 2370
box -8 -3 16 105
use FILL  FILL_564
timestamp 1714281807
transform 1 0 2984 0 1 2370
box -8 -3 16 105
use FILL  FILL_565
timestamp 1714281807
transform 1 0 2976 0 1 2370
box -8 -3 16 105
use FILL  FILL_566
timestamp 1714281807
transform 1 0 2968 0 1 2370
box -8 -3 16 105
use FILL  FILL_567
timestamp 1714281807
transform 1 0 2960 0 1 2370
box -8 -3 16 105
use FILL  FILL_568
timestamp 1714281807
transform 1 0 2952 0 1 2370
box -8 -3 16 105
use FILL  FILL_569
timestamp 1714281807
transform 1 0 2944 0 1 2370
box -8 -3 16 105
use FILL  FILL_570
timestamp 1714281807
transform 1 0 2936 0 1 2370
box -8 -3 16 105
use FILL  FILL_571
timestamp 1714281807
transform 1 0 2928 0 1 2370
box -8 -3 16 105
use FILL  FILL_572
timestamp 1714281807
transform 1 0 2920 0 1 2370
box -8 -3 16 105
use FILL  FILL_573
timestamp 1714281807
transform 1 0 2912 0 1 2370
box -8 -3 16 105
use FILL  FILL_574
timestamp 1714281807
transform 1 0 2808 0 1 2370
box -8 -3 16 105
use FILL  FILL_575
timestamp 1714281807
transform 1 0 2800 0 1 2370
box -8 -3 16 105
use FILL  FILL_576
timestamp 1714281807
transform 1 0 2792 0 1 2370
box -8 -3 16 105
use FILL  FILL_577
timestamp 1714281807
transform 1 0 2760 0 1 2370
box -8 -3 16 105
use FILL  FILL_578
timestamp 1714281807
transform 1 0 2752 0 1 2370
box -8 -3 16 105
use FILL  FILL_579
timestamp 1714281807
transform 1 0 2744 0 1 2370
box -8 -3 16 105
use FILL  FILL_580
timestamp 1714281807
transform 1 0 2736 0 1 2370
box -8 -3 16 105
use FILL  FILL_581
timestamp 1714281807
transform 1 0 2728 0 1 2370
box -8 -3 16 105
use FILL  FILL_582
timestamp 1714281807
transform 1 0 2720 0 1 2370
box -8 -3 16 105
use FILL  FILL_583
timestamp 1714281807
transform 1 0 2680 0 1 2370
box -8 -3 16 105
use FILL  FILL_584
timestamp 1714281807
transform 1 0 2672 0 1 2370
box -8 -3 16 105
use FILL  FILL_585
timestamp 1714281807
transform 1 0 2664 0 1 2370
box -8 -3 16 105
use FILL  FILL_586
timestamp 1714281807
transform 1 0 2640 0 1 2370
box -8 -3 16 105
use FILL  FILL_587
timestamp 1714281807
transform 1 0 2632 0 1 2370
box -8 -3 16 105
use FILL  FILL_588
timestamp 1714281807
transform 1 0 2624 0 1 2370
box -8 -3 16 105
use FILL  FILL_589
timestamp 1714281807
transform 1 0 2584 0 1 2370
box -8 -3 16 105
use FILL  FILL_590
timestamp 1714281807
transform 1 0 2576 0 1 2370
box -8 -3 16 105
use FILL  FILL_591
timestamp 1714281807
transform 1 0 2568 0 1 2370
box -8 -3 16 105
use FILL  FILL_592
timestamp 1714281807
transform 1 0 2560 0 1 2370
box -8 -3 16 105
use FILL  FILL_593
timestamp 1714281807
transform 1 0 2552 0 1 2370
box -8 -3 16 105
use FILL  FILL_594
timestamp 1714281807
transform 1 0 2544 0 1 2370
box -8 -3 16 105
use FILL  FILL_595
timestamp 1714281807
transform 1 0 2512 0 1 2370
box -8 -3 16 105
use FILL  FILL_596
timestamp 1714281807
transform 1 0 2504 0 1 2370
box -8 -3 16 105
use FILL  FILL_597
timestamp 1714281807
transform 1 0 2496 0 1 2370
box -8 -3 16 105
use FILL  FILL_598
timestamp 1714281807
transform 1 0 2456 0 1 2370
box -8 -3 16 105
use FILL  FILL_599
timestamp 1714281807
transform 1 0 2448 0 1 2370
box -8 -3 16 105
use FILL  FILL_600
timestamp 1714281807
transform 1 0 2440 0 1 2370
box -8 -3 16 105
use FILL  FILL_601
timestamp 1714281807
transform 1 0 2432 0 1 2370
box -8 -3 16 105
use FILL  FILL_602
timestamp 1714281807
transform 1 0 2424 0 1 2370
box -8 -3 16 105
use FILL  FILL_603
timestamp 1714281807
transform 1 0 2416 0 1 2370
box -8 -3 16 105
use FILL  FILL_604
timestamp 1714281807
transform 1 0 2384 0 1 2370
box -8 -3 16 105
use FILL  FILL_605
timestamp 1714281807
transform 1 0 2376 0 1 2370
box -8 -3 16 105
use FILL  FILL_606
timestamp 1714281807
transform 1 0 2368 0 1 2370
box -8 -3 16 105
use FILL  FILL_607
timestamp 1714281807
transform 1 0 2360 0 1 2370
box -8 -3 16 105
use FILL  FILL_608
timestamp 1714281807
transform 1 0 2320 0 1 2370
box -8 -3 16 105
use FILL  FILL_609
timestamp 1714281807
transform 1 0 2312 0 1 2370
box -8 -3 16 105
use FILL  FILL_610
timestamp 1714281807
transform 1 0 2304 0 1 2370
box -8 -3 16 105
use FILL  FILL_611
timestamp 1714281807
transform 1 0 2296 0 1 2370
box -8 -3 16 105
use FILL  FILL_612
timestamp 1714281807
transform 1 0 2288 0 1 2370
box -8 -3 16 105
use FILL  FILL_613
timestamp 1714281807
transform 1 0 2256 0 1 2370
box -8 -3 16 105
use FILL  FILL_614
timestamp 1714281807
transform 1 0 2248 0 1 2370
box -8 -3 16 105
use FILL  FILL_615
timestamp 1714281807
transform 1 0 2240 0 1 2370
box -8 -3 16 105
use FILL  FILL_616
timestamp 1714281807
transform 1 0 2232 0 1 2370
box -8 -3 16 105
use FILL  FILL_617
timestamp 1714281807
transform 1 0 2192 0 1 2370
box -8 -3 16 105
use FILL  FILL_618
timestamp 1714281807
transform 1 0 2184 0 1 2370
box -8 -3 16 105
use FILL  FILL_619
timestamp 1714281807
transform 1 0 2176 0 1 2370
box -8 -3 16 105
use FILL  FILL_620
timestamp 1714281807
transform 1 0 2168 0 1 2370
box -8 -3 16 105
use FILL  FILL_621
timestamp 1714281807
transform 1 0 2160 0 1 2370
box -8 -3 16 105
use FILL  FILL_622
timestamp 1714281807
transform 1 0 2152 0 1 2370
box -8 -3 16 105
use FILL  FILL_623
timestamp 1714281807
transform 1 0 2144 0 1 2370
box -8 -3 16 105
use FILL  FILL_624
timestamp 1714281807
transform 1 0 2088 0 1 2370
box -8 -3 16 105
use FILL  FILL_625
timestamp 1714281807
transform 1 0 2080 0 1 2370
box -8 -3 16 105
use FILL  FILL_626
timestamp 1714281807
transform 1 0 2072 0 1 2370
box -8 -3 16 105
use FILL  FILL_627
timestamp 1714281807
transform 1 0 2064 0 1 2370
box -8 -3 16 105
use FILL  FILL_628
timestamp 1714281807
transform 1 0 2056 0 1 2370
box -8 -3 16 105
use FILL  FILL_629
timestamp 1714281807
transform 1 0 2048 0 1 2370
box -8 -3 16 105
use FILL  FILL_630
timestamp 1714281807
transform 1 0 2040 0 1 2370
box -8 -3 16 105
use FILL  FILL_631
timestamp 1714281807
transform 1 0 2008 0 1 2370
box -8 -3 16 105
use FILL  FILL_632
timestamp 1714281807
transform 1 0 2000 0 1 2370
box -8 -3 16 105
use FILL  FILL_633
timestamp 1714281807
transform 1 0 1992 0 1 2370
box -8 -3 16 105
use FILL  FILL_634
timestamp 1714281807
transform 1 0 1984 0 1 2370
box -8 -3 16 105
use FILL  FILL_635
timestamp 1714281807
transform 1 0 1944 0 1 2370
box -8 -3 16 105
use FILL  FILL_636
timestamp 1714281807
transform 1 0 1936 0 1 2370
box -8 -3 16 105
use FILL  FILL_637
timestamp 1714281807
transform 1 0 1928 0 1 2370
box -8 -3 16 105
use FILL  FILL_638
timestamp 1714281807
transform 1 0 1824 0 1 2370
box -8 -3 16 105
use FILL  FILL_639
timestamp 1714281807
transform 1 0 1816 0 1 2370
box -8 -3 16 105
use FILL  FILL_640
timestamp 1714281807
transform 1 0 1808 0 1 2370
box -8 -3 16 105
use FILL  FILL_641
timestamp 1714281807
transform 1 0 1768 0 1 2370
box -8 -3 16 105
use FILL  FILL_642
timestamp 1714281807
transform 1 0 1760 0 1 2370
box -8 -3 16 105
use FILL  FILL_643
timestamp 1714281807
transform 1 0 1728 0 1 2370
box -8 -3 16 105
use FILL  FILL_644
timestamp 1714281807
transform 1 0 1720 0 1 2370
box -8 -3 16 105
use FILL  FILL_645
timestamp 1714281807
transform 1 0 1712 0 1 2370
box -8 -3 16 105
use FILL  FILL_646
timestamp 1714281807
transform 1 0 1704 0 1 2370
box -8 -3 16 105
use FILL  FILL_647
timestamp 1714281807
transform 1 0 1600 0 1 2370
box -8 -3 16 105
use FILL  FILL_648
timestamp 1714281807
transform 1 0 1592 0 1 2370
box -8 -3 16 105
use FILL  FILL_649
timestamp 1714281807
transform 1 0 1584 0 1 2370
box -8 -3 16 105
use FILL  FILL_650
timestamp 1714281807
transform 1 0 1552 0 1 2370
box -8 -3 16 105
use FILL  FILL_651
timestamp 1714281807
transform 1 0 1544 0 1 2370
box -8 -3 16 105
use FILL  FILL_652
timestamp 1714281807
transform 1 0 1536 0 1 2370
box -8 -3 16 105
use FILL  FILL_653
timestamp 1714281807
transform 1 0 1528 0 1 2370
box -8 -3 16 105
use FILL  FILL_654
timestamp 1714281807
transform 1 0 1488 0 1 2370
box -8 -3 16 105
use FILL  FILL_655
timestamp 1714281807
transform 1 0 1480 0 1 2370
box -8 -3 16 105
use FILL  FILL_656
timestamp 1714281807
transform 1 0 1472 0 1 2370
box -8 -3 16 105
use FILL  FILL_657
timestamp 1714281807
transform 1 0 1464 0 1 2370
box -8 -3 16 105
use FILL  FILL_658
timestamp 1714281807
transform 1 0 1456 0 1 2370
box -8 -3 16 105
use FILL  FILL_659
timestamp 1714281807
transform 1 0 1448 0 1 2370
box -8 -3 16 105
use FILL  FILL_660
timestamp 1714281807
transform 1 0 1408 0 1 2370
box -8 -3 16 105
use FILL  FILL_661
timestamp 1714281807
transform 1 0 1400 0 1 2370
box -8 -3 16 105
use FILL  FILL_662
timestamp 1714281807
transform 1 0 1392 0 1 2370
box -8 -3 16 105
use FILL  FILL_663
timestamp 1714281807
transform 1 0 1384 0 1 2370
box -8 -3 16 105
use FILL  FILL_664
timestamp 1714281807
transform 1 0 1280 0 1 2370
box -8 -3 16 105
use FILL  FILL_665
timestamp 1714281807
transform 1 0 1272 0 1 2370
box -8 -3 16 105
use FILL  FILL_666
timestamp 1714281807
transform 1 0 1168 0 1 2370
box -8 -3 16 105
use FILL  FILL_667
timestamp 1714281807
transform 1 0 1160 0 1 2370
box -8 -3 16 105
use FILL  FILL_668
timestamp 1714281807
transform 1 0 1056 0 1 2370
box -8 -3 16 105
use FILL  FILL_669
timestamp 1714281807
transform 1 0 952 0 1 2370
box -8 -3 16 105
use FILL  FILL_670
timestamp 1714281807
transform 1 0 944 0 1 2370
box -8 -3 16 105
use FILL  FILL_671
timestamp 1714281807
transform 1 0 936 0 1 2370
box -8 -3 16 105
use FILL  FILL_672
timestamp 1714281807
transform 1 0 904 0 1 2370
box -8 -3 16 105
use FILL  FILL_673
timestamp 1714281807
transform 1 0 896 0 1 2370
box -8 -3 16 105
use FILL  FILL_674
timestamp 1714281807
transform 1 0 888 0 1 2370
box -8 -3 16 105
use FILL  FILL_675
timestamp 1714281807
transform 1 0 880 0 1 2370
box -8 -3 16 105
use FILL  FILL_676
timestamp 1714281807
transform 1 0 872 0 1 2370
box -8 -3 16 105
use FILL  FILL_677
timestamp 1714281807
transform 1 0 840 0 1 2370
box -8 -3 16 105
use FILL  FILL_678
timestamp 1714281807
transform 1 0 832 0 1 2370
box -8 -3 16 105
use FILL  FILL_679
timestamp 1714281807
transform 1 0 824 0 1 2370
box -8 -3 16 105
use FILL  FILL_680
timestamp 1714281807
transform 1 0 816 0 1 2370
box -8 -3 16 105
use FILL  FILL_681
timestamp 1714281807
transform 1 0 808 0 1 2370
box -8 -3 16 105
use FILL  FILL_682
timestamp 1714281807
transform 1 0 800 0 1 2370
box -8 -3 16 105
use FILL  FILL_683
timestamp 1714281807
transform 1 0 768 0 1 2370
box -8 -3 16 105
use FILL  FILL_684
timestamp 1714281807
transform 1 0 760 0 1 2370
box -8 -3 16 105
use FILL  FILL_685
timestamp 1714281807
transform 1 0 752 0 1 2370
box -8 -3 16 105
use FILL  FILL_686
timestamp 1714281807
transform 1 0 744 0 1 2370
box -8 -3 16 105
use FILL  FILL_687
timestamp 1714281807
transform 1 0 736 0 1 2370
box -8 -3 16 105
use FILL  FILL_688
timestamp 1714281807
transform 1 0 696 0 1 2370
box -8 -3 16 105
use FILL  FILL_689
timestamp 1714281807
transform 1 0 688 0 1 2370
box -8 -3 16 105
use FILL  FILL_690
timestamp 1714281807
transform 1 0 680 0 1 2370
box -8 -3 16 105
use FILL  FILL_691
timestamp 1714281807
transform 1 0 656 0 1 2370
box -8 -3 16 105
use FILL  FILL_692
timestamp 1714281807
transform 1 0 648 0 1 2370
box -8 -3 16 105
use FILL  FILL_693
timestamp 1714281807
transform 1 0 544 0 1 2370
box -8 -3 16 105
use FILL  FILL_694
timestamp 1714281807
transform 1 0 536 0 1 2370
box -8 -3 16 105
use FILL  FILL_695
timestamp 1714281807
transform 1 0 528 0 1 2370
box -8 -3 16 105
use FILL  FILL_696
timestamp 1714281807
transform 1 0 520 0 1 2370
box -8 -3 16 105
use FILL  FILL_697
timestamp 1714281807
transform 1 0 488 0 1 2370
box -8 -3 16 105
use FILL  FILL_698
timestamp 1714281807
transform 1 0 480 0 1 2370
box -8 -3 16 105
use FILL  FILL_699
timestamp 1714281807
transform 1 0 472 0 1 2370
box -8 -3 16 105
use FILL  FILL_700
timestamp 1714281807
transform 1 0 464 0 1 2370
box -8 -3 16 105
use FILL  FILL_701
timestamp 1714281807
transform 1 0 456 0 1 2370
box -8 -3 16 105
use FILL  FILL_702
timestamp 1714281807
transform 1 0 448 0 1 2370
box -8 -3 16 105
use FILL  FILL_703
timestamp 1714281807
transform 1 0 416 0 1 2370
box -8 -3 16 105
use FILL  FILL_704
timestamp 1714281807
transform 1 0 408 0 1 2370
box -8 -3 16 105
use FILL  FILL_705
timestamp 1714281807
transform 1 0 400 0 1 2370
box -8 -3 16 105
use FILL  FILL_706
timestamp 1714281807
transform 1 0 392 0 1 2370
box -8 -3 16 105
use FILL  FILL_707
timestamp 1714281807
transform 1 0 384 0 1 2370
box -8 -3 16 105
use FILL  FILL_708
timestamp 1714281807
transform 1 0 376 0 1 2370
box -8 -3 16 105
use FILL  FILL_709
timestamp 1714281807
transform 1 0 344 0 1 2370
box -8 -3 16 105
use FILL  FILL_710
timestamp 1714281807
transform 1 0 336 0 1 2370
box -8 -3 16 105
use FILL  FILL_711
timestamp 1714281807
transform 1 0 328 0 1 2370
box -8 -3 16 105
use FILL  FILL_712
timestamp 1714281807
transform 1 0 320 0 1 2370
box -8 -3 16 105
use FILL  FILL_713
timestamp 1714281807
transform 1 0 312 0 1 2370
box -8 -3 16 105
use FILL  FILL_714
timestamp 1714281807
transform 1 0 304 0 1 2370
box -8 -3 16 105
use FILL  FILL_715
timestamp 1714281807
transform 1 0 296 0 1 2370
box -8 -3 16 105
use FILL  FILL_716
timestamp 1714281807
transform 1 0 248 0 1 2370
box -8 -3 16 105
use FILL  FILL_717
timestamp 1714281807
transform 1 0 240 0 1 2370
box -8 -3 16 105
use FILL  FILL_718
timestamp 1714281807
transform 1 0 232 0 1 2370
box -8 -3 16 105
use FILL  FILL_719
timestamp 1714281807
transform 1 0 224 0 1 2370
box -8 -3 16 105
use FILL  FILL_720
timestamp 1714281807
transform 1 0 216 0 1 2370
box -8 -3 16 105
use FILL  FILL_721
timestamp 1714281807
transform 1 0 208 0 1 2370
box -8 -3 16 105
use FILL  FILL_722
timestamp 1714281807
transform 1 0 200 0 1 2370
box -8 -3 16 105
use FILL  FILL_723
timestamp 1714281807
transform 1 0 192 0 1 2370
box -8 -3 16 105
use FILL  FILL_724
timestamp 1714281807
transform 1 0 184 0 1 2370
box -8 -3 16 105
use FILL  FILL_725
timestamp 1714281807
transform 1 0 176 0 1 2370
box -8 -3 16 105
use FILL  FILL_726
timestamp 1714281807
transform 1 0 168 0 1 2370
box -8 -3 16 105
use FILL  FILL_727
timestamp 1714281807
transform 1 0 160 0 1 2370
box -8 -3 16 105
use FILL  FILL_728
timestamp 1714281807
transform 1 0 152 0 1 2370
box -8 -3 16 105
use FILL  FILL_729
timestamp 1714281807
transform 1 0 144 0 1 2370
box -8 -3 16 105
use FILL  FILL_730
timestamp 1714281807
transform 1 0 136 0 1 2370
box -8 -3 16 105
use FILL  FILL_731
timestamp 1714281807
transform 1 0 128 0 1 2370
box -8 -3 16 105
use FILL  FILL_732
timestamp 1714281807
transform 1 0 120 0 1 2370
box -8 -3 16 105
use FILL  FILL_733
timestamp 1714281807
transform 1 0 112 0 1 2370
box -8 -3 16 105
use FILL  FILL_734
timestamp 1714281807
transform 1 0 104 0 1 2370
box -8 -3 16 105
use FILL  FILL_735
timestamp 1714281807
transform 1 0 96 0 1 2370
box -8 -3 16 105
use FILL  FILL_736
timestamp 1714281807
transform 1 0 88 0 1 2370
box -8 -3 16 105
use FILL  FILL_737
timestamp 1714281807
transform 1 0 80 0 1 2370
box -8 -3 16 105
use FILL  FILL_738
timestamp 1714281807
transform 1 0 72 0 1 2370
box -8 -3 16 105
use FILL  FILL_739
timestamp 1714281807
transform 1 0 3000 0 -1 2370
box -8 -3 16 105
use FILL  FILL_740
timestamp 1714281807
transform 1 0 2992 0 -1 2370
box -8 -3 16 105
use FILL  FILL_741
timestamp 1714281807
transform 1 0 2984 0 -1 2370
box -8 -3 16 105
use FILL  FILL_742
timestamp 1714281807
transform 1 0 2976 0 -1 2370
box -8 -3 16 105
use FILL  FILL_743
timestamp 1714281807
transform 1 0 2968 0 -1 2370
box -8 -3 16 105
use FILL  FILL_744
timestamp 1714281807
transform 1 0 2960 0 -1 2370
box -8 -3 16 105
use FILL  FILL_745
timestamp 1714281807
transform 1 0 2952 0 -1 2370
box -8 -3 16 105
use FILL  FILL_746
timestamp 1714281807
transform 1 0 2944 0 -1 2370
box -8 -3 16 105
use FILL  FILL_747
timestamp 1714281807
transform 1 0 2936 0 -1 2370
box -8 -3 16 105
use FILL  FILL_748
timestamp 1714281807
transform 1 0 2928 0 -1 2370
box -8 -3 16 105
use FILL  FILL_749
timestamp 1714281807
transform 1 0 2920 0 -1 2370
box -8 -3 16 105
use FILL  FILL_750
timestamp 1714281807
transform 1 0 2912 0 -1 2370
box -8 -3 16 105
use FILL  FILL_751
timestamp 1714281807
transform 1 0 2904 0 -1 2370
box -8 -3 16 105
use FILL  FILL_752
timestamp 1714281807
transform 1 0 2896 0 -1 2370
box -8 -3 16 105
use FILL  FILL_753
timestamp 1714281807
transform 1 0 2888 0 -1 2370
box -8 -3 16 105
use FILL  FILL_754
timestamp 1714281807
transform 1 0 2880 0 -1 2370
box -8 -3 16 105
use FILL  FILL_755
timestamp 1714281807
transform 1 0 2872 0 -1 2370
box -8 -3 16 105
use FILL  FILL_756
timestamp 1714281807
transform 1 0 2864 0 -1 2370
box -8 -3 16 105
use FILL  FILL_757
timestamp 1714281807
transform 1 0 2760 0 -1 2370
box -8 -3 16 105
use FILL  FILL_758
timestamp 1714281807
transform 1 0 2752 0 -1 2370
box -8 -3 16 105
use FILL  FILL_759
timestamp 1714281807
transform 1 0 2728 0 -1 2370
box -8 -3 16 105
use FILL  FILL_760
timestamp 1714281807
transform 1 0 2720 0 -1 2370
box -8 -3 16 105
use FILL  FILL_761
timestamp 1714281807
transform 1 0 2712 0 -1 2370
box -8 -3 16 105
use FILL  FILL_762
timestamp 1714281807
transform 1 0 2704 0 -1 2370
box -8 -3 16 105
use FILL  FILL_763
timestamp 1714281807
transform 1 0 2672 0 -1 2370
box -8 -3 16 105
use FILL  FILL_764
timestamp 1714281807
transform 1 0 2664 0 -1 2370
box -8 -3 16 105
use FILL  FILL_765
timestamp 1714281807
transform 1 0 2560 0 -1 2370
box -8 -3 16 105
use FILL  FILL_766
timestamp 1714281807
transform 1 0 2456 0 -1 2370
box -8 -3 16 105
use FILL  FILL_767
timestamp 1714281807
transform 1 0 2448 0 -1 2370
box -8 -3 16 105
use FILL  FILL_768
timestamp 1714281807
transform 1 0 2440 0 -1 2370
box -8 -3 16 105
use FILL  FILL_769
timestamp 1714281807
transform 1 0 2336 0 -1 2370
box -8 -3 16 105
use FILL  FILL_770
timestamp 1714281807
transform 1 0 2328 0 -1 2370
box -8 -3 16 105
use FILL  FILL_771
timestamp 1714281807
transform 1 0 2224 0 -1 2370
box -8 -3 16 105
use FILL  FILL_772
timestamp 1714281807
transform 1 0 2216 0 -1 2370
box -8 -3 16 105
use FILL  FILL_773
timestamp 1714281807
transform 1 0 2208 0 -1 2370
box -8 -3 16 105
use FILL  FILL_774
timestamp 1714281807
transform 1 0 2200 0 -1 2370
box -8 -3 16 105
use FILL  FILL_775
timestamp 1714281807
transform 1 0 2192 0 -1 2370
box -8 -3 16 105
use FILL  FILL_776
timestamp 1714281807
transform 1 0 2184 0 -1 2370
box -8 -3 16 105
use FILL  FILL_777
timestamp 1714281807
transform 1 0 2176 0 -1 2370
box -8 -3 16 105
use FILL  FILL_778
timestamp 1714281807
transform 1 0 2168 0 -1 2370
box -8 -3 16 105
use FILL  FILL_779
timestamp 1714281807
transform 1 0 2160 0 -1 2370
box -8 -3 16 105
use FILL  FILL_780
timestamp 1714281807
transform 1 0 2104 0 -1 2370
box -8 -3 16 105
use FILL  FILL_781
timestamp 1714281807
transform 1 0 2096 0 -1 2370
box -8 -3 16 105
use FILL  FILL_782
timestamp 1714281807
transform 1 0 2088 0 -1 2370
box -8 -3 16 105
use FILL  FILL_783
timestamp 1714281807
transform 1 0 1984 0 -1 2370
box -8 -3 16 105
use FILL  FILL_784
timestamp 1714281807
transform 1 0 1976 0 -1 2370
box -8 -3 16 105
use FILL  FILL_785
timestamp 1714281807
transform 1 0 1944 0 -1 2370
box -8 -3 16 105
use FILL  FILL_786
timestamp 1714281807
transform 1 0 1936 0 -1 2370
box -8 -3 16 105
use FILL  FILL_787
timestamp 1714281807
transform 1 0 1928 0 -1 2370
box -8 -3 16 105
use FILL  FILL_788
timestamp 1714281807
transform 1 0 1920 0 -1 2370
box -8 -3 16 105
use FILL  FILL_789
timestamp 1714281807
transform 1 0 1912 0 -1 2370
box -8 -3 16 105
use FILL  FILL_790
timestamp 1714281807
transform 1 0 1904 0 -1 2370
box -8 -3 16 105
use FILL  FILL_791
timestamp 1714281807
transform 1 0 1848 0 -1 2370
box -8 -3 16 105
use FILL  FILL_792
timestamp 1714281807
transform 1 0 1840 0 -1 2370
box -8 -3 16 105
use FILL  FILL_793
timestamp 1714281807
transform 1 0 1616 0 -1 2370
box -8 -3 16 105
use FILL  FILL_794
timestamp 1714281807
transform 1 0 1608 0 -1 2370
box -8 -3 16 105
use FILL  FILL_795
timestamp 1714281807
transform 1 0 1600 0 -1 2370
box -8 -3 16 105
use FILL  FILL_796
timestamp 1714281807
transform 1 0 1592 0 -1 2370
box -8 -3 16 105
use FILL  FILL_797
timestamp 1714281807
transform 1 0 1536 0 -1 2370
box -8 -3 16 105
use FILL  FILL_798
timestamp 1714281807
transform 1 0 1528 0 -1 2370
box -8 -3 16 105
use FILL  FILL_799
timestamp 1714281807
transform 1 0 1424 0 -1 2370
box -8 -3 16 105
use FILL  FILL_800
timestamp 1714281807
transform 1 0 1416 0 -1 2370
box -8 -3 16 105
use FILL  FILL_801
timestamp 1714281807
transform 1 0 1408 0 -1 2370
box -8 -3 16 105
use FILL  FILL_802
timestamp 1714281807
transform 1 0 1352 0 -1 2370
box -8 -3 16 105
use FILL  FILL_803
timestamp 1714281807
transform 1 0 1344 0 -1 2370
box -8 -3 16 105
use FILL  FILL_804
timestamp 1714281807
transform 1 0 1336 0 -1 2370
box -8 -3 16 105
use FILL  FILL_805
timestamp 1714281807
transform 1 0 1328 0 -1 2370
box -8 -3 16 105
use FILL  FILL_806
timestamp 1714281807
transform 1 0 1320 0 -1 2370
box -8 -3 16 105
use FILL  FILL_807
timestamp 1714281807
transform 1 0 1312 0 -1 2370
box -8 -3 16 105
use FILL  FILL_808
timestamp 1714281807
transform 1 0 1256 0 -1 2370
box -8 -3 16 105
use FILL  FILL_809
timestamp 1714281807
transform 1 0 1248 0 -1 2370
box -8 -3 16 105
use FILL  FILL_810
timestamp 1714281807
transform 1 0 1240 0 -1 2370
box -8 -3 16 105
use FILL  FILL_811
timestamp 1714281807
transform 1 0 1232 0 -1 2370
box -8 -3 16 105
use FILL  FILL_812
timestamp 1714281807
transform 1 0 1224 0 -1 2370
box -8 -3 16 105
use FILL  FILL_813
timestamp 1714281807
transform 1 0 1216 0 -1 2370
box -8 -3 16 105
use FILL  FILL_814
timestamp 1714281807
transform 1 0 1208 0 -1 2370
box -8 -3 16 105
use FILL  FILL_815
timestamp 1714281807
transform 1 0 1200 0 -1 2370
box -8 -3 16 105
use FILL  FILL_816
timestamp 1714281807
transform 1 0 1192 0 -1 2370
box -8 -3 16 105
use FILL  FILL_817
timestamp 1714281807
transform 1 0 1136 0 -1 2370
box -8 -3 16 105
use FILL  FILL_818
timestamp 1714281807
transform 1 0 1128 0 -1 2370
box -8 -3 16 105
use FILL  FILL_819
timestamp 1714281807
transform 1 0 1120 0 -1 2370
box -8 -3 16 105
use FILL  FILL_820
timestamp 1714281807
transform 1 0 1112 0 -1 2370
box -8 -3 16 105
use FILL  FILL_821
timestamp 1714281807
transform 1 0 1088 0 -1 2370
box -8 -3 16 105
use FILL  FILL_822
timestamp 1714281807
transform 1 0 1080 0 -1 2370
box -8 -3 16 105
use FILL  FILL_823
timestamp 1714281807
transform 1 0 1040 0 -1 2370
box -8 -3 16 105
use FILL  FILL_824
timestamp 1714281807
transform 1 0 1032 0 -1 2370
box -8 -3 16 105
use FILL  FILL_825
timestamp 1714281807
transform 1 0 1024 0 -1 2370
box -8 -3 16 105
use FILL  FILL_826
timestamp 1714281807
transform 1 0 1016 0 -1 2370
box -8 -3 16 105
use FILL  FILL_827
timestamp 1714281807
transform 1 0 1008 0 -1 2370
box -8 -3 16 105
use FILL  FILL_828
timestamp 1714281807
transform 1 0 1000 0 -1 2370
box -8 -3 16 105
use FILL  FILL_829
timestamp 1714281807
transform 1 0 992 0 -1 2370
box -8 -3 16 105
use FILL  FILL_830
timestamp 1714281807
transform 1 0 952 0 -1 2370
box -8 -3 16 105
use FILL  FILL_831
timestamp 1714281807
transform 1 0 944 0 -1 2370
box -8 -3 16 105
use FILL  FILL_832
timestamp 1714281807
transform 1 0 936 0 -1 2370
box -8 -3 16 105
use FILL  FILL_833
timestamp 1714281807
transform 1 0 928 0 -1 2370
box -8 -3 16 105
use FILL  FILL_834
timestamp 1714281807
transform 1 0 920 0 -1 2370
box -8 -3 16 105
use FILL  FILL_835
timestamp 1714281807
transform 1 0 816 0 -1 2370
box -8 -3 16 105
use FILL  FILL_836
timestamp 1714281807
transform 1 0 808 0 -1 2370
box -8 -3 16 105
use FILL  FILL_837
timestamp 1714281807
transform 1 0 704 0 -1 2370
box -8 -3 16 105
use FILL  FILL_838
timestamp 1714281807
transform 1 0 600 0 -1 2370
box -8 -3 16 105
use FILL  FILL_839
timestamp 1714281807
transform 1 0 496 0 -1 2370
box -8 -3 16 105
use FILL  FILL_840
timestamp 1714281807
transform 1 0 488 0 -1 2370
box -8 -3 16 105
use FILL  FILL_841
timestamp 1714281807
transform 1 0 480 0 -1 2370
box -8 -3 16 105
use FILL  FILL_842
timestamp 1714281807
transform 1 0 448 0 -1 2370
box -8 -3 16 105
use FILL  FILL_843
timestamp 1714281807
transform 1 0 440 0 -1 2370
box -8 -3 16 105
use FILL  FILL_844
timestamp 1714281807
transform 1 0 432 0 -1 2370
box -8 -3 16 105
use FILL  FILL_845
timestamp 1714281807
transform 1 0 408 0 -1 2370
box -8 -3 16 105
use FILL  FILL_846
timestamp 1714281807
transform 1 0 400 0 -1 2370
box -8 -3 16 105
use FILL  FILL_847
timestamp 1714281807
transform 1 0 392 0 -1 2370
box -8 -3 16 105
use FILL  FILL_848
timestamp 1714281807
transform 1 0 384 0 -1 2370
box -8 -3 16 105
use FILL  FILL_849
timestamp 1714281807
transform 1 0 376 0 -1 2370
box -8 -3 16 105
use FILL  FILL_850
timestamp 1714281807
transform 1 0 344 0 -1 2370
box -8 -3 16 105
use FILL  FILL_851
timestamp 1714281807
transform 1 0 336 0 -1 2370
box -8 -3 16 105
use FILL  FILL_852
timestamp 1714281807
transform 1 0 328 0 -1 2370
box -8 -3 16 105
use FILL  FILL_853
timestamp 1714281807
transform 1 0 320 0 -1 2370
box -8 -3 16 105
use FILL  FILL_854
timestamp 1714281807
transform 1 0 312 0 -1 2370
box -8 -3 16 105
use FILL  FILL_855
timestamp 1714281807
transform 1 0 304 0 -1 2370
box -8 -3 16 105
use FILL  FILL_856
timestamp 1714281807
transform 1 0 280 0 -1 2370
box -8 -3 16 105
use FILL  FILL_857
timestamp 1714281807
transform 1 0 272 0 -1 2370
box -8 -3 16 105
use FILL  FILL_858
timestamp 1714281807
transform 1 0 168 0 -1 2370
box -8 -3 16 105
use FILL  FILL_859
timestamp 1714281807
transform 1 0 160 0 -1 2370
box -8 -3 16 105
use FILL  FILL_860
timestamp 1714281807
transform 1 0 152 0 -1 2370
box -8 -3 16 105
use FILL  FILL_861
timestamp 1714281807
transform 1 0 144 0 -1 2370
box -8 -3 16 105
use FILL  FILL_862
timestamp 1714281807
transform 1 0 136 0 -1 2370
box -8 -3 16 105
use FILL  FILL_863
timestamp 1714281807
transform 1 0 128 0 -1 2370
box -8 -3 16 105
use FILL  FILL_864
timestamp 1714281807
transform 1 0 120 0 -1 2370
box -8 -3 16 105
use FILL  FILL_865
timestamp 1714281807
transform 1 0 112 0 -1 2370
box -8 -3 16 105
use FILL  FILL_866
timestamp 1714281807
transform 1 0 104 0 -1 2370
box -8 -3 16 105
use FILL  FILL_867
timestamp 1714281807
transform 1 0 96 0 -1 2370
box -8 -3 16 105
use FILL  FILL_868
timestamp 1714281807
transform 1 0 88 0 -1 2370
box -8 -3 16 105
use FILL  FILL_869
timestamp 1714281807
transform 1 0 80 0 -1 2370
box -8 -3 16 105
use FILL  FILL_870
timestamp 1714281807
transform 1 0 72 0 -1 2370
box -8 -3 16 105
use FILL  FILL_871
timestamp 1714281807
transform 1 0 3000 0 1 2170
box -8 -3 16 105
use FILL  FILL_872
timestamp 1714281807
transform 1 0 2992 0 1 2170
box -8 -3 16 105
use FILL  FILL_873
timestamp 1714281807
transform 1 0 2984 0 1 2170
box -8 -3 16 105
use FILL  FILL_874
timestamp 1714281807
transform 1 0 2976 0 1 2170
box -8 -3 16 105
use FILL  FILL_875
timestamp 1714281807
transform 1 0 2968 0 1 2170
box -8 -3 16 105
use FILL  FILL_876
timestamp 1714281807
transform 1 0 2960 0 1 2170
box -8 -3 16 105
use FILL  FILL_877
timestamp 1714281807
transform 1 0 2952 0 1 2170
box -8 -3 16 105
use FILL  FILL_878
timestamp 1714281807
transform 1 0 2848 0 1 2170
box -8 -3 16 105
use FILL  FILL_879
timestamp 1714281807
transform 1 0 2840 0 1 2170
box -8 -3 16 105
use FILL  FILL_880
timestamp 1714281807
transform 1 0 2816 0 1 2170
box -8 -3 16 105
use FILL  FILL_881
timestamp 1714281807
transform 1 0 2808 0 1 2170
box -8 -3 16 105
use FILL  FILL_882
timestamp 1714281807
transform 1 0 2800 0 1 2170
box -8 -3 16 105
use FILL  FILL_883
timestamp 1714281807
transform 1 0 2792 0 1 2170
box -8 -3 16 105
use FILL  FILL_884
timestamp 1714281807
transform 1 0 2784 0 1 2170
box -8 -3 16 105
use FILL  FILL_885
timestamp 1714281807
transform 1 0 2744 0 1 2170
box -8 -3 16 105
use FILL  FILL_886
timestamp 1714281807
transform 1 0 2736 0 1 2170
box -8 -3 16 105
use FILL  FILL_887
timestamp 1714281807
transform 1 0 2728 0 1 2170
box -8 -3 16 105
use FILL  FILL_888
timestamp 1714281807
transform 1 0 2664 0 1 2170
box -8 -3 16 105
use FILL  FILL_889
timestamp 1714281807
transform 1 0 2656 0 1 2170
box -8 -3 16 105
use FILL  FILL_890
timestamp 1714281807
transform 1 0 2624 0 1 2170
box -8 -3 16 105
use FILL  FILL_891
timestamp 1714281807
transform 1 0 2616 0 1 2170
box -8 -3 16 105
use FILL  FILL_892
timestamp 1714281807
transform 1 0 2608 0 1 2170
box -8 -3 16 105
use FILL  FILL_893
timestamp 1714281807
transform 1 0 2504 0 1 2170
box -8 -3 16 105
use FILL  FILL_894
timestamp 1714281807
transform 1 0 2400 0 1 2170
box -8 -3 16 105
use FILL  FILL_895
timestamp 1714281807
transform 1 0 2392 0 1 2170
box -8 -3 16 105
use FILL  FILL_896
timestamp 1714281807
transform 1 0 2384 0 1 2170
box -8 -3 16 105
use FILL  FILL_897
timestamp 1714281807
transform 1 0 2344 0 1 2170
box -8 -3 16 105
use FILL  FILL_898
timestamp 1714281807
transform 1 0 2336 0 1 2170
box -8 -3 16 105
use FILL  FILL_899
timestamp 1714281807
transform 1 0 2328 0 1 2170
box -8 -3 16 105
use FILL  FILL_900
timestamp 1714281807
transform 1 0 2320 0 1 2170
box -8 -3 16 105
use FILL  FILL_901
timestamp 1714281807
transform 1 0 2312 0 1 2170
box -8 -3 16 105
use FILL  FILL_902
timestamp 1714281807
transform 1 0 2280 0 1 2170
box -8 -3 16 105
use FILL  FILL_903
timestamp 1714281807
transform 1 0 2272 0 1 2170
box -8 -3 16 105
use FILL  FILL_904
timestamp 1714281807
transform 1 0 2264 0 1 2170
box -8 -3 16 105
use FILL  FILL_905
timestamp 1714281807
transform 1 0 2256 0 1 2170
box -8 -3 16 105
use FILL  FILL_906
timestamp 1714281807
transform 1 0 2248 0 1 2170
box -8 -3 16 105
use FILL  FILL_907
timestamp 1714281807
transform 1 0 2240 0 1 2170
box -8 -3 16 105
use FILL  FILL_908
timestamp 1714281807
transform 1 0 2232 0 1 2170
box -8 -3 16 105
use FILL  FILL_909
timestamp 1714281807
transform 1 0 2192 0 1 2170
box -8 -3 16 105
use FILL  FILL_910
timestamp 1714281807
transform 1 0 2184 0 1 2170
box -8 -3 16 105
use FILL  FILL_911
timestamp 1714281807
transform 1 0 2176 0 1 2170
box -8 -3 16 105
use FILL  FILL_912
timestamp 1714281807
transform 1 0 2168 0 1 2170
box -8 -3 16 105
use FILL  FILL_913
timestamp 1714281807
transform 1 0 2064 0 1 2170
box -8 -3 16 105
use FILL  FILL_914
timestamp 1714281807
transform 1 0 2056 0 1 2170
box -8 -3 16 105
use FILL  FILL_915
timestamp 1714281807
transform 1 0 2048 0 1 2170
box -8 -3 16 105
use FILL  FILL_916
timestamp 1714281807
transform 1 0 2040 0 1 2170
box -8 -3 16 105
use FILL  FILL_917
timestamp 1714281807
transform 1 0 2016 0 1 2170
box -8 -3 16 105
use FILL  FILL_918
timestamp 1714281807
transform 1 0 2008 0 1 2170
box -8 -3 16 105
use FILL  FILL_919
timestamp 1714281807
transform 1 0 2000 0 1 2170
box -8 -3 16 105
use FILL  FILL_920
timestamp 1714281807
transform 1 0 1936 0 1 2170
box -8 -3 16 105
use FILL  FILL_921
timestamp 1714281807
transform 1 0 1928 0 1 2170
box -8 -3 16 105
use FILL  FILL_922
timestamp 1714281807
transform 1 0 1920 0 1 2170
box -8 -3 16 105
use FILL  FILL_923
timestamp 1714281807
transform 1 0 1856 0 1 2170
box -8 -3 16 105
use FILL  FILL_924
timestamp 1714281807
transform 1 0 1848 0 1 2170
box -8 -3 16 105
use FILL  FILL_925
timestamp 1714281807
transform 1 0 1840 0 1 2170
box -8 -3 16 105
use FILL  FILL_926
timestamp 1714281807
transform 1 0 1800 0 1 2170
box -8 -3 16 105
use FILL  FILL_927
timestamp 1714281807
transform 1 0 1792 0 1 2170
box -8 -3 16 105
use FILL  FILL_928
timestamp 1714281807
transform 1 0 1784 0 1 2170
box -8 -3 16 105
use FILL  FILL_929
timestamp 1714281807
transform 1 0 1776 0 1 2170
box -8 -3 16 105
use FILL  FILL_930
timestamp 1714281807
transform 1 0 1768 0 1 2170
box -8 -3 16 105
use FILL  FILL_931
timestamp 1714281807
transform 1 0 1760 0 1 2170
box -8 -3 16 105
use FILL  FILL_932
timestamp 1714281807
transform 1 0 1752 0 1 2170
box -8 -3 16 105
use FILL  FILL_933
timestamp 1714281807
transform 1 0 1728 0 1 2170
box -8 -3 16 105
use FILL  FILL_934
timestamp 1714281807
transform 1 0 1720 0 1 2170
box -8 -3 16 105
use FILL  FILL_935
timestamp 1714281807
transform 1 0 1696 0 1 2170
box -8 -3 16 105
use FILL  FILL_936
timestamp 1714281807
transform 1 0 1688 0 1 2170
box -8 -3 16 105
use FILL  FILL_937
timestamp 1714281807
transform 1 0 1680 0 1 2170
box -8 -3 16 105
use FILL  FILL_938
timestamp 1714281807
transform 1 0 1672 0 1 2170
box -8 -3 16 105
use FILL  FILL_939
timestamp 1714281807
transform 1 0 1664 0 1 2170
box -8 -3 16 105
use FILL  FILL_940
timestamp 1714281807
transform 1 0 1656 0 1 2170
box -8 -3 16 105
use FILL  FILL_941
timestamp 1714281807
transform 1 0 1648 0 1 2170
box -8 -3 16 105
use FILL  FILL_942
timestamp 1714281807
transform 1 0 1616 0 1 2170
box -8 -3 16 105
use FILL  FILL_943
timestamp 1714281807
transform 1 0 1608 0 1 2170
box -8 -3 16 105
use FILL  FILL_944
timestamp 1714281807
transform 1 0 1600 0 1 2170
box -8 -3 16 105
use FILL  FILL_945
timestamp 1714281807
transform 1 0 1592 0 1 2170
box -8 -3 16 105
use FILL  FILL_946
timestamp 1714281807
transform 1 0 1584 0 1 2170
box -8 -3 16 105
use FILL  FILL_947
timestamp 1714281807
transform 1 0 1576 0 1 2170
box -8 -3 16 105
use FILL  FILL_948
timestamp 1714281807
transform 1 0 1568 0 1 2170
box -8 -3 16 105
use FILL  FILL_949
timestamp 1714281807
transform 1 0 1560 0 1 2170
box -8 -3 16 105
use FILL  FILL_950
timestamp 1714281807
transform 1 0 1496 0 1 2170
box -8 -3 16 105
use FILL  FILL_951
timestamp 1714281807
transform 1 0 1488 0 1 2170
box -8 -3 16 105
use FILL  FILL_952
timestamp 1714281807
transform 1 0 1480 0 1 2170
box -8 -3 16 105
use FILL  FILL_953
timestamp 1714281807
transform 1 0 1376 0 1 2170
box -8 -3 16 105
use FILL  FILL_954
timestamp 1714281807
transform 1 0 1368 0 1 2170
box -8 -3 16 105
use FILL  FILL_955
timestamp 1714281807
transform 1 0 1360 0 1 2170
box -8 -3 16 105
use FILL  FILL_956
timestamp 1714281807
transform 1 0 1336 0 1 2170
box -8 -3 16 105
use FILL  FILL_957
timestamp 1714281807
transform 1 0 1328 0 1 2170
box -8 -3 16 105
use FILL  FILL_958
timestamp 1714281807
transform 1 0 1320 0 1 2170
box -8 -3 16 105
use FILL  FILL_959
timestamp 1714281807
transform 1 0 1312 0 1 2170
box -8 -3 16 105
use FILL  FILL_960
timestamp 1714281807
transform 1 0 1304 0 1 2170
box -8 -3 16 105
use FILL  FILL_961
timestamp 1714281807
transform 1 0 1256 0 1 2170
box -8 -3 16 105
use FILL  FILL_962
timestamp 1714281807
transform 1 0 1248 0 1 2170
box -8 -3 16 105
use FILL  FILL_963
timestamp 1714281807
transform 1 0 1240 0 1 2170
box -8 -3 16 105
use FILL  FILL_964
timestamp 1714281807
transform 1 0 1232 0 1 2170
box -8 -3 16 105
use FILL  FILL_965
timestamp 1714281807
transform 1 0 1224 0 1 2170
box -8 -3 16 105
use FILL  FILL_966
timestamp 1714281807
transform 1 0 1216 0 1 2170
box -8 -3 16 105
use FILL  FILL_967
timestamp 1714281807
transform 1 0 1176 0 1 2170
box -8 -3 16 105
use FILL  FILL_968
timestamp 1714281807
transform 1 0 1168 0 1 2170
box -8 -3 16 105
use FILL  FILL_969
timestamp 1714281807
transform 1 0 1160 0 1 2170
box -8 -3 16 105
use FILL  FILL_970
timestamp 1714281807
transform 1 0 1152 0 1 2170
box -8 -3 16 105
use FILL  FILL_971
timestamp 1714281807
transform 1 0 1144 0 1 2170
box -8 -3 16 105
use FILL  FILL_972
timestamp 1714281807
transform 1 0 1104 0 1 2170
box -8 -3 16 105
use FILL  FILL_973
timestamp 1714281807
transform 1 0 1096 0 1 2170
box -8 -3 16 105
use FILL  FILL_974
timestamp 1714281807
transform 1 0 1088 0 1 2170
box -8 -3 16 105
use FILL  FILL_975
timestamp 1714281807
transform 1 0 1080 0 1 2170
box -8 -3 16 105
use FILL  FILL_976
timestamp 1714281807
transform 1 0 1072 0 1 2170
box -8 -3 16 105
use FILL  FILL_977
timestamp 1714281807
transform 1 0 1064 0 1 2170
box -8 -3 16 105
use FILL  FILL_978
timestamp 1714281807
transform 1 0 1032 0 1 2170
box -8 -3 16 105
use FILL  FILL_979
timestamp 1714281807
transform 1 0 1024 0 1 2170
box -8 -3 16 105
use FILL  FILL_980
timestamp 1714281807
transform 1 0 1016 0 1 2170
box -8 -3 16 105
use FILL  FILL_981
timestamp 1714281807
transform 1 0 976 0 1 2170
box -8 -3 16 105
use FILL  FILL_982
timestamp 1714281807
transform 1 0 968 0 1 2170
box -8 -3 16 105
use FILL  FILL_983
timestamp 1714281807
transform 1 0 960 0 1 2170
box -8 -3 16 105
use FILL  FILL_984
timestamp 1714281807
transform 1 0 952 0 1 2170
box -8 -3 16 105
use FILL  FILL_985
timestamp 1714281807
transform 1 0 944 0 1 2170
box -8 -3 16 105
use FILL  FILL_986
timestamp 1714281807
transform 1 0 936 0 1 2170
box -8 -3 16 105
use FILL  FILL_987
timestamp 1714281807
transform 1 0 928 0 1 2170
box -8 -3 16 105
use FILL  FILL_988
timestamp 1714281807
transform 1 0 888 0 1 2170
box -8 -3 16 105
use FILL  FILL_989
timestamp 1714281807
transform 1 0 880 0 1 2170
box -8 -3 16 105
use FILL  FILL_990
timestamp 1714281807
transform 1 0 872 0 1 2170
box -8 -3 16 105
use FILL  FILL_991
timestamp 1714281807
transform 1 0 864 0 1 2170
box -8 -3 16 105
use FILL  FILL_992
timestamp 1714281807
transform 1 0 856 0 1 2170
box -8 -3 16 105
use FILL  FILL_993
timestamp 1714281807
transform 1 0 832 0 1 2170
box -8 -3 16 105
use FILL  FILL_994
timestamp 1714281807
transform 1 0 728 0 1 2170
box -8 -3 16 105
use FILL  FILL_995
timestamp 1714281807
transform 1 0 704 0 1 2170
box -8 -3 16 105
use FILL  FILL_996
timestamp 1714281807
transform 1 0 696 0 1 2170
box -8 -3 16 105
use FILL  FILL_997
timestamp 1714281807
transform 1 0 688 0 1 2170
box -8 -3 16 105
use FILL  FILL_998
timestamp 1714281807
transform 1 0 584 0 1 2170
box -8 -3 16 105
use FILL  FILL_999
timestamp 1714281807
transform 1 0 576 0 1 2170
box -8 -3 16 105
use FILL  FILL_1000
timestamp 1714281807
transform 1 0 472 0 1 2170
box -8 -3 16 105
use FILL  FILL_1001
timestamp 1714281807
transform 1 0 464 0 1 2170
box -8 -3 16 105
use FILL  FILL_1002
timestamp 1714281807
transform 1 0 456 0 1 2170
box -8 -3 16 105
use FILL  FILL_1003
timestamp 1714281807
transform 1 0 448 0 1 2170
box -8 -3 16 105
use FILL  FILL_1004
timestamp 1714281807
transform 1 0 408 0 1 2170
box -8 -3 16 105
use FILL  FILL_1005
timestamp 1714281807
transform 1 0 384 0 1 2170
box -8 -3 16 105
use FILL  FILL_1006
timestamp 1714281807
transform 1 0 376 0 1 2170
box -8 -3 16 105
use FILL  FILL_1007
timestamp 1714281807
transform 1 0 368 0 1 2170
box -8 -3 16 105
use FILL  FILL_1008
timestamp 1714281807
transform 1 0 360 0 1 2170
box -8 -3 16 105
use FILL  FILL_1009
timestamp 1714281807
transform 1 0 256 0 1 2170
box -8 -3 16 105
use FILL  FILL_1010
timestamp 1714281807
transform 1 0 248 0 1 2170
box -8 -3 16 105
use FILL  FILL_1011
timestamp 1714281807
transform 1 0 240 0 1 2170
box -8 -3 16 105
use FILL  FILL_1012
timestamp 1714281807
transform 1 0 232 0 1 2170
box -8 -3 16 105
use FILL  FILL_1013
timestamp 1714281807
transform 1 0 224 0 1 2170
box -8 -3 16 105
use FILL  FILL_1014
timestamp 1714281807
transform 1 0 216 0 1 2170
box -8 -3 16 105
use FILL  FILL_1015
timestamp 1714281807
transform 1 0 208 0 1 2170
box -8 -3 16 105
use FILL  FILL_1016
timestamp 1714281807
transform 1 0 200 0 1 2170
box -8 -3 16 105
use FILL  FILL_1017
timestamp 1714281807
transform 1 0 192 0 1 2170
box -8 -3 16 105
use FILL  FILL_1018
timestamp 1714281807
transform 1 0 184 0 1 2170
box -8 -3 16 105
use FILL  FILL_1019
timestamp 1714281807
transform 1 0 176 0 1 2170
box -8 -3 16 105
use FILL  FILL_1020
timestamp 1714281807
transform 1 0 168 0 1 2170
box -8 -3 16 105
use FILL  FILL_1021
timestamp 1714281807
transform 1 0 160 0 1 2170
box -8 -3 16 105
use FILL  FILL_1022
timestamp 1714281807
transform 1 0 152 0 1 2170
box -8 -3 16 105
use FILL  FILL_1023
timestamp 1714281807
transform 1 0 144 0 1 2170
box -8 -3 16 105
use FILL  FILL_1024
timestamp 1714281807
transform 1 0 136 0 1 2170
box -8 -3 16 105
use FILL  FILL_1025
timestamp 1714281807
transform 1 0 128 0 1 2170
box -8 -3 16 105
use FILL  FILL_1026
timestamp 1714281807
transform 1 0 120 0 1 2170
box -8 -3 16 105
use FILL  FILL_1027
timestamp 1714281807
transform 1 0 112 0 1 2170
box -8 -3 16 105
use FILL  FILL_1028
timestamp 1714281807
transform 1 0 104 0 1 2170
box -8 -3 16 105
use FILL  FILL_1029
timestamp 1714281807
transform 1 0 96 0 1 2170
box -8 -3 16 105
use FILL  FILL_1030
timestamp 1714281807
transform 1 0 88 0 1 2170
box -8 -3 16 105
use FILL  FILL_1031
timestamp 1714281807
transform 1 0 80 0 1 2170
box -8 -3 16 105
use FILL  FILL_1032
timestamp 1714281807
transform 1 0 72 0 1 2170
box -8 -3 16 105
use FILL  FILL_1033
timestamp 1714281807
transform 1 0 3000 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1034
timestamp 1714281807
transform 1 0 2992 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1035
timestamp 1714281807
transform 1 0 2984 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1036
timestamp 1714281807
transform 1 0 2976 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1037
timestamp 1714281807
transform 1 0 2968 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1038
timestamp 1714281807
transform 1 0 2960 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1039
timestamp 1714281807
transform 1 0 2952 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1040
timestamp 1714281807
transform 1 0 2944 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1041
timestamp 1714281807
transform 1 0 2936 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1042
timestamp 1714281807
transform 1 0 2928 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1043
timestamp 1714281807
transform 1 0 2920 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1044
timestamp 1714281807
transform 1 0 2912 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1045
timestamp 1714281807
transform 1 0 2872 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1046
timestamp 1714281807
transform 1 0 2864 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1047
timestamp 1714281807
transform 1 0 2856 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1048
timestamp 1714281807
transform 1 0 2848 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1049
timestamp 1714281807
transform 1 0 2840 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1050
timestamp 1714281807
transform 1 0 2792 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1051
timestamp 1714281807
transform 1 0 2784 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1052
timestamp 1714281807
transform 1 0 2776 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1053
timestamp 1714281807
transform 1 0 2768 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1054
timestamp 1714281807
transform 1 0 2760 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1055
timestamp 1714281807
transform 1 0 2712 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1056
timestamp 1714281807
transform 1 0 2704 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1057
timestamp 1714281807
transform 1 0 2696 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1058
timestamp 1714281807
transform 1 0 2688 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1059
timestamp 1714281807
transform 1 0 2592 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1060
timestamp 1714281807
transform 1 0 2584 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1061
timestamp 1714281807
transform 1 0 2576 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1062
timestamp 1714281807
transform 1 0 2472 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1063
timestamp 1714281807
transform 1 0 2464 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1064
timestamp 1714281807
transform 1 0 2456 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1065
timestamp 1714281807
transform 1 0 2408 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1066
timestamp 1714281807
transform 1 0 2400 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1067
timestamp 1714281807
transform 1 0 2392 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1068
timestamp 1714281807
transform 1 0 2384 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1069
timestamp 1714281807
transform 1 0 2320 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1070
timestamp 1714281807
transform 1 0 2312 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1071
timestamp 1714281807
transform 1 0 2272 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1072
timestamp 1714281807
transform 1 0 2264 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1073
timestamp 1714281807
transform 1 0 2256 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1074
timestamp 1714281807
transform 1 0 2248 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1075
timestamp 1714281807
transform 1 0 2224 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1076
timestamp 1714281807
transform 1 0 2216 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1077
timestamp 1714281807
transform 1 0 2112 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1078
timestamp 1714281807
transform 1 0 2080 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1079
timestamp 1714281807
transform 1 0 2072 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1080
timestamp 1714281807
transform 1 0 2064 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1081
timestamp 1714281807
transform 1 0 2056 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1082
timestamp 1714281807
transform 1 0 2048 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1083
timestamp 1714281807
transform 1 0 2000 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1084
timestamp 1714281807
transform 1 0 1992 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1085
timestamp 1714281807
transform 1 0 1984 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1086
timestamp 1714281807
transform 1 0 1976 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1087
timestamp 1714281807
transform 1 0 1968 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1088
timestamp 1714281807
transform 1 0 1920 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1089
timestamp 1714281807
transform 1 0 1912 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1090
timestamp 1714281807
transform 1 0 1904 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1091
timestamp 1714281807
transform 1 0 1896 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1092
timestamp 1714281807
transform 1 0 1888 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1093
timestamp 1714281807
transform 1 0 1864 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1094
timestamp 1714281807
transform 1 0 1824 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1095
timestamp 1714281807
transform 1 0 1816 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1096
timestamp 1714281807
transform 1 0 1808 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1097
timestamp 1714281807
transform 1 0 1800 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1098
timestamp 1714281807
transform 1 0 1792 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1099
timestamp 1714281807
transform 1 0 1760 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1100
timestamp 1714281807
transform 1 0 1752 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1101
timestamp 1714281807
transform 1 0 1712 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1102
timestamp 1714281807
transform 1 0 1704 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1103
timestamp 1714281807
transform 1 0 1696 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1104
timestamp 1714281807
transform 1 0 1688 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1105
timestamp 1714281807
transform 1 0 1680 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1106
timestamp 1714281807
transform 1 0 1672 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1107
timestamp 1714281807
transform 1 0 1616 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1108
timestamp 1714281807
transform 1 0 1608 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1109
timestamp 1714281807
transform 1 0 1600 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1110
timestamp 1714281807
transform 1 0 1592 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1111
timestamp 1714281807
transform 1 0 1584 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1112
timestamp 1714281807
transform 1 0 1552 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1113
timestamp 1714281807
transform 1 0 1544 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1114
timestamp 1714281807
transform 1 0 1536 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1115
timestamp 1714281807
transform 1 0 1496 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1116
timestamp 1714281807
transform 1 0 1488 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1117
timestamp 1714281807
transform 1 0 1480 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1118
timestamp 1714281807
transform 1 0 1472 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1119
timestamp 1714281807
transform 1 0 1368 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1120
timestamp 1714281807
transform 1 0 1360 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1121
timestamp 1714281807
transform 1 0 1336 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1122
timestamp 1714281807
transform 1 0 1328 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1123
timestamp 1714281807
transform 1 0 1320 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1124
timestamp 1714281807
transform 1 0 1312 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1125
timestamp 1714281807
transform 1 0 1264 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1126
timestamp 1714281807
transform 1 0 1256 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1127
timestamp 1714281807
transform 1 0 1248 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1128
timestamp 1714281807
transform 1 0 1240 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1129
timestamp 1714281807
transform 1 0 1232 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1130
timestamp 1714281807
transform 1 0 1200 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1131
timestamp 1714281807
transform 1 0 1192 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1132
timestamp 1714281807
transform 1 0 1152 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1133
timestamp 1714281807
transform 1 0 1144 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1134
timestamp 1714281807
transform 1 0 1040 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1135
timestamp 1714281807
transform 1 0 1032 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1136
timestamp 1714281807
transform 1 0 992 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1137
timestamp 1714281807
transform 1 0 984 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1138
timestamp 1714281807
transform 1 0 944 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1139
timestamp 1714281807
transform 1 0 936 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1140
timestamp 1714281807
transform 1 0 928 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1141
timestamp 1714281807
transform 1 0 888 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1142
timestamp 1714281807
transform 1 0 880 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1143
timestamp 1714281807
transform 1 0 872 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1144
timestamp 1714281807
transform 1 0 864 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1145
timestamp 1714281807
transform 1 0 856 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1146
timestamp 1714281807
transform 1 0 816 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1147
timestamp 1714281807
transform 1 0 808 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1148
timestamp 1714281807
transform 1 0 784 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1149
timestamp 1714281807
transform 1 0 776 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1150
timestamp 1714281807
transform 1 0 768 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1151
timestamp 1714281807
transform 1 0 760 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1152
timestamp 1714281807
transform 1 0 752 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1153
timestamp 1714281807
transform 1 0 712 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1154
timestamp 1714281807
transform 1 0 704 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1155
timestamp 1714281807
transform 1 0 696 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1156
timestamp 1714281807
transform 1 0 664 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1157
timestamp 1714281807
transform 1 0 656 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1158
timestamp 1714281807
transform 1 0 648 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1159
timestamp 1714281807
transform 1 0 640 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1160
timestamp 1714281807
transform 1 0 632 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1161
timestamp 1714281807
transform 1 0 624 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1162
timestamp 1714281807
transform 1 0 584 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1163
timestamp 1714281807
transform 1 0 576 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1164
timestamp 1714281807
transform 1 0 552 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1165
timestamp 1714281807
transform 1 0 544 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1166
timestamp 1714281807
transform 1 0 536 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1167
timestamp 1714281807
transform 1 0 528 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1168
timestamp 1714281807
transform 1 0 520 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1169
timestamp 1714281807
transform 1 0 488 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1170
timestamp 1714281807
transform 1 0 480 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1171
timestamp 1714281807
transform 1 0 472 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1172
timestamp 1714281807
transform 1 0 464 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1173
timestamp 1714281807
transform 1 0 424 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1174
timestamp 1714281807
transform 1 0 416 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1175
timestamp 1714281807
transform 1 0 408 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1176
timestamp 1714281807
transform 1 0 304 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1177
timestamp 1714281807
transform 1 0 296 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1178
timestamp 1714281807
transform 1 0 192 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1179
timestamp 1714281807
transform 1 0 184 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1180
timestamp 1714281807
transform 1 0 176 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1181
timestamp 1714281807
transform 1 0 168 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1182
timestamp 1714281807
transform 1 0 160 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1183
timestamp 1714281807
transform 1 0 152 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1184
timestamp 1714281807
transform 1 0 144 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1185
timestamp 1714281807
transform 1 0 136 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1186
timestamp 1714281807
transform 1 0 128 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1187
timestamp 1714281807
transform 1 0 120 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1188
timestamp 1714281807
transform 1 0 112 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1189
timestamp 1714281807
transform 1 0 104 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1190
timestamp 1714281807
transform 1 0 96 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1191
timestamp 1714281807
transform 1 0 88 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1192
timestamp 1714281807
transform 1 0 80 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1193
timestamp 1714281807
transform 1 0 72 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1194
timestamp 1714281807
transform 1 0 3000 0 1 1970
box -8 -3 16 105
use FILL  FILL_1195
timestamp 1714281807
transform 1 0 2896 0 1 1970
box -8 -3 16 105
use FILL  FILL_1196
timestamp 1714281807
transform 1 0 2888 0 1 1970
box -8 -3 16 105
use FILL  FILL_1197
timestamp 1714281807
transform 1 0 2832 0 1 1970
box -8 -3 16 105
use FILL  FILL_1198
timestamp 1714281807
transform 1 0 2824 0 1 1970
box -8 -3 16 105
use FILL  FILL_1199
timestamp 1714281807
transform 1 0 2816 0 1 1970
box -8 -3 16 105
use FILL  FILL_1200
timestamp 1714281807
transform 1 0 2808 0 1 1970
box -8 -3 16 105
use FILL  FILL_1201
timestamp 1714281807
transform 1 0 2800 0 1 1970
box -8 -3 16 105
use FILL  FILL_1202
timestamp 1714281807
transform 1 0 2792 0 1 1970
box -8 -3 16 105
use FILL  FILL_1203
timestamp 1714281807
transform 1 0 2784 0 1 1970
box -8 -3 16 105
use FILL  FILL_1204
timestamp 1714281807
transform 1 0 2736 0 1 1970
box -8 -3 16 105
use FILL  FILL_1205
timestamp 1714281807
transform 1 0 2728 0 1 1970
box -8 -3 16 105
use FILL  FILL_1206
timestamp 1714281807
transform 1 0 2720 0 1 1970
box -8 -3 16 105
use FILL  FILL_1207
timestamp 1714281807
transform 1 0 2712 0 1 1970
box -8 -3 16 105
use FILL  FILL_1208
timestamp 1714281807
transform 1 0 2616 0 1 1970
box -8 -3 16 105
use FILL  FILL_1209
timestamp 1714281807
transform 1 0 2608 0 1 1970
box -8 -3 16 105
use FILL  FILL_1210
timestamp 1714281807
transform 1 0 2576 0 1 1970
box -8 -3 16 105
use FILL  FILL_1211
timestamp 1714281807
transform 1 0 2568 0 1 1970
box -8 -3 16 105
use FILL  FILL_1212
timestamp 1714281807
transform 1 0 2464 0 1 1970
box -8 -3 16 105
use FILL  FILL_1213
timestamp 1714281807
transform 1 0 2456 0 1 1970
box -8 -3 16 105
use FILL  FILL_1214
timestamp 1714281807
transform 1 0 2448 0 1 1970
box -8 -3 16 105
use FILL  FILL_1215
timestamp 1714281807
transform 1 0 2408 0 1 1970
box -8 -3 16 105
use FILL  FILL_1216
timestamp 1714281807
transform 1 0 2400 0 1 1970
box -8 -3 16 105
use FILL  FILL_1217
timestamp 1714281807
transform 1 0 2392 0 1 1970
box -8 -3 16 105
use FILL  FILL_1218
timestamp 1714281807
transform 1 0 2384 0 1 1970
box -8 -3 16 105
use FILL  FILL_1219
timestamp 1714281807
transform 1 0 2376 0 1 1970
box -8 -3 16 105
use FILL  FILL_1220
timestamp 1714281807
transform 1 0 2368 0 1 1970
box -8 -3 16 105
use FILL  FILL_1221
timestamp 1714281807
transform 1 0 2360 0 1 1970
box -8 -3 16 105
use FILL  FILL_1222
timestamp 1714281807
transform 1 0 2312 0 1 1970
box -8 -3 16 105
use FILL  FILL_1223
timestamp 1714281807
transform 1 0 2304 0 1 1970
box -8 -3 16 105
use FILL  FILL_1224
timestamp 1714281807
transform 1 0 2296 0 1 1970
box -8 -3 16 105
use FILL  FILL_1225
timestamp 1714281807
transform 1 0 2288 0 1 1970
box -8 -3 16 105
use FILL  FILL_1226
timestamp 1714281807
transform 1 0 2184 0 1 1970
box -8 -3 16 105
use FILL  FILL_1227
timestamp 1714281807
transform 1 0 2176 0 1 1970
box -8 -3 16 105
use FILL  FILL_1228
timestamp 1714281807
transform 1 0 2168 0 1 1970
box -8 -3 16 105
use FILL  FILL_1229
timestamp 1714281807
transform 1 0 2160 0 1 1970
box -8 -3 16 105
use FILL  FILL_1230
timestamp 1714281807
transform 1 0 2120 0 1 1970
box -8 -3 16 105
use FILL  FILL_1231
timestamp 1714281807
transform 1 0 2112 0 1 1970
box -8 -3 16 105
use FILL  FILL_1232
timestamp 1714281807
transform 1 0 2104 0 1 1970
box -8 -3 16 105
use FILL  FILL_1233
timestamp 1714281807
transform 1 0 2096 0 1 1970
box -8 -3 16 105
use FILL  FILL_1234
timestamp 1714281807
transform 1 0 2088 0 1 1970
box -8 -3 16 105
use FILL  FILL_1235
timestamp 1714281807
transform 1 0 2080 0 1 1970
box -8 -3 16 105
use FILL  FILL_1236
timestamp 1714281807
transform 1 0 2072 0 1 1970
box -8 -3 16 105
use FILL  FILL_1237
timestamp 1714281807
transform 1 0 2024 0 1 1970
box -8 -3 16 105
use FILL  FILL_1238
timestamp 1714281807
transform 1 0 2016 0 1 1970
box -8 -3 16 105
use FILL  FILL_1239
timestamp 1714281807
transform 1 0 2008 0 1 1970
box -8 -3 16 105
use FILL  FILL_1240
timestamp 1714281807
transform 1 0 2000 0 1 1970
box -8 -3 16 105
use FILL  FILL_1241
timestamp 1714281807
transform 1 0 1992 0 1 1970
box -8 -3 16 105
use FILL  FILL_1242
timestamp 1714281807
transform 1 0 1984 0 1 1970
box -8 -3 16 105
use FILL  FILL_1243
timestamp 1714281807
transform 1 0 1976 0 1 1970
box -8 -3 16 105
use FILL  FILL_1244
timestamp 1714281807
transform 1 0 1928 0 1 1970
box -8 -3 16 105
use FILL  FILL_1245
timestamp 1714281807
transform 1 0 1920 0 1 1970
box -8 -3 16 105
use FILL  FILL_1246
timestamp 1714281807
transform 1 0 1912 0 1 1970
box -8 -3 16 105
use FILL  FILL_1247
timestamp 1714281807
transform 1 0 1888 0 1 1970
box -8 -3 16 105
use FILL  FILL_1248
timestamp 1714281807
transform 1 0 1880 0 1 1970
box -8 -3 16 105
use FILL  FILL_1249
timestamp 1714281807
transform 1 0 1872 0 1 1970
box -8 -3 16 105
use FILL  FILL_1250
timestamp 1714281807
transform 1 0 1864 0 1 1970
box -8 -3 16 105
use FILL  FILL_1251
timestamp 1714281807
transform 1 0 1824 0 1 1970
box -8 -3 16 105
use FILL  FILL_1252
timestamp 1714281807
transform 1 0 1816 0 1 1970
box -8 -3 16 105
use FILL  FILL_1253
timestamp 1714281807
transform 1 0 1776 0 1 1970
box -8 -3 16 105
use FILL  FILL_1254
timestamp 1714281807
transform 1 0 1768 0 1 1970
box -8 -3 16 105
use FILL  FILL_1255
timestamp 1714281807
transform 1 0 1760 0 1 1970
box -8 -3 16 105
use FILL  FILL_1256
timestamp 1714281807
transform 1 0 1752 0 1 1970
box -8 -3 16 105
use FILL  FILL_1257
timestamp 1714281807
transform 1 0 1744 0 1 1970
box -8 -3 16 105
use FILL  FILL_1258
timestamp 1714281807
transform 1 0 1736 0 1 1970
box -8 -3 16 105
use FILL  FILL_1259
timestamp 1714281807
transform 1 0 1728 0 1 1970
box -8 -3 16 105
use FILL  FILL_1260
timestamp 1714281807
transform 1 0 1680 0 1 1970
box -8 -3 16 105
use FILL  FILL_1261
timestamp 1714281807
transform 1 0 1672 0 1 1970
box -8 -3 16 105
use FILL  FILL_1262
timestamp 1714281807
transform 1 0 1664 0 1 1970
box -8 -3 16 105
use FILL  FILL_1263
timestamp 1714281807
transform 1 0 1656 0 1 1970
box -8 -3 16 105
use FILL  FILL_1264
timestamp 1714281807
transform 1 0 1648 0 1 1970
box -8 -3 16 105
use FILL  FILL_1265
timestamp 1714281807
transform 1 0 1640 0 1 1970
box -8 -3 16 105
use FILL  FILL_1266
timestamp 1714281807
transform 1 0 1560 0 1 1970
box -8 -3 16 105
use FILL  FILL_1267
timestamp 1714281807
transform 1 0 1552 0 1 1970
box -8 -3 16 105
use FILL  FILL_1268
timestamp 1714281807
transform 1 0 1544 0 1 1970
box -8 -3 16 105
use FILL  FILL_1269
timestamp 1714281807
transform 1 0 1512 0 1 1970
box -8 -3 16 105
use FILL  FILL_1270
timestamp 1714281807
transform 1 0 1504 0 1 1970
box -8 -3 16 105
use FILL  FILL_1271
timestamp 1714281807
transform 1 0 1496 0 1 1970
box -8 -3 16 105
use FILL  FILL_1272
timestamp 1714281807
transform 1 0 1488 0 1 1970
box -8 -3 16 105
use FILL  FILL_1273
timestamp 1714281807
transform 1 0 1456 0 1 1970
box -8 -3 16 105
use FILL  FILL_1274
timestamp 1714281807
transform 1 0 1448 0 1 1970
box -8 -3 16 105
use FILL  FILL_1275
timestamp 1714281807
transform 1 0 1440 0 1 1970
box -8 -3 16 105
use FILL  FILL_1276
timestamp 1714281807
transform 1 0 1432 0 1 1970
box -8 -3 16 105
use FILL  FILL_1277
timestamp 1714281807
transform 1 0 1408 0 1 1970
box -8 -3 16 105
use FILL  FILL_1278
timestamp 1714281807
transform 1 0 1400 0 1 1970
box -8 -3 16 105
use FILL  FILL_1279
timestamp 1714281807
transform 1 0 1392 0 1 1970
box -8 -3 16 105
use FILL  FILL_1280
timestamp 1714281807
transform 1 0 1344 0 1 1970
box -8 -3 16 105
use FILL  FILL_1281
timestamp 1714281807
transform 1 0 1336 0 1 1970
box -8 -3 16 105
use FILL  FILL_1282
timestamp 1714281807
transform 1 0 1328 0 1 1970
box -8 -3 16 105
use FILL  FILL_1283
timestamp 1714281807
transform 1 0 1320 0 1 1970
box -8 -3 16 105
use FILL  FILL_1284
timestamp 1714281807
transform 1 0 1312 0 1 1970
box -8 -3 16 105
use FILL  FILL_1285
timestamp 1714281807
transform 1 0 1304 0 1 1970
box -8 -3 16 105
use FILL  FILL_1286
timestamp 1714281807
transform 1 0 1256 0 1 1970
box -8 -3 16 105
use FILL  FILL_1287
timestamp 1714281807
transform 1 0 1248 0 1 1970
box -8 -3 16 105
use FILL  FILL_1288
timestamp 1714281807
transform 1 0 1240 0 1 1970
box -8 -3 16 105
use FILL  FILL_1289
timestamp 1714281807
transform 1 0 1216 0 1 1970
box -8 -3 16 105
use FILL  FILL_1290
timestamp 1714281807
transform 1 0 1208 0 1 1970
box -8 -3 16 105
use FILL  FILL_1291
timestamp 1714281807
transform 1 0 1200 0 1 1970
box -8 -3 16 105
use FILL  FILL_1292
timestamp 1714281807
transform 1 0 1168 0 1 1970
box -8 -3 16 105
use FILL  FILL_1293
timestamp 1714281807
transform 1 0 1160 0 1 1970
box -8 -3 16 105
use FILL  FILL_1294
timestamp 1714281807
transform 1 0 1120 0 1 1970
box -8 -3 16 105
use FILL  FILL_1295
timestamp 1714281807
transform 1 0 1112 0 1 1970
box -8 -3 16 105
use FILL  FILL_1296
timestamp 1714281807
transform 1 0 1008 0 1 1970
box -8 -3 16 105
use FILL  FILL_1297
timestamp 1714281807
transform 1 0 984 0 1 1970
box -8 -3 16 105
use FILL  FILL_1298
timestamp 1714281807
transform 1 0 976 0 1 1970
box -8 -3 16 105
use FILL  FILL_1299
timestamp 1714281807
transform 1 0 928 0 1 1970
box -8 -3 16 105
use FILL  FILL_1300
timestamp 1714281807
transform 1 0 920 0 1 1970
box -8 -3 16 105
use FILL  FILL_1301
timestamp 1714281807
transform 1 0 792 0 1 1970
box -8 -3 16 105
use FILL  FILL_1302
timestamp 1714281807
transform 1 0 784 0 1 1970
box -8 -3 16 105
use FILL  FILL_1303
timestamp 1714281807
transform 1 0 680 0 1 1970
box -8 -3 16 105
use FILL  FILL_1304
timestamp 1714281807
transform 1 0 672 0 1 1970
box -8 -3 16 105
use FILL  FILL_1305
timestamp 1714281807
transform 1 0 664 0 1 1970
box -8 -3 16 105
use FILL  FILL_1306
timestamp 1714281807
transform 1 0 656 0 1 1970
box -8 -3 16 105
use FILL  FILL_1307
timestamp 1714281807
transform 1 0 616 0 1 1970
box -8 -3 16 105
use FILL  FILL_1308
timestamp 1714281807
transform 1 0 592 0 1 1970
box -8 -3 16 105
use FILL  FILL_1309
timestamp 1714281807
transform 1 0 584 0 1 1970
box -8 -3 16 105
use FILL  FILL_1310
timestamp 1714281807
transform 1 0 576 0 1 1970
box -8 -3 16 105
use FILL  FILL_1311
timestamp 1714281807
transform 1 0 568 0 1 1970
box -8 -3 16 105
use FILL  FILL_1312
timestamp 1714281807
transform 1 0 528 0 1 1970
box -8 -3 16 105
use FILL  FILL_1313
timestamp 1714281807
transform 1 0 520 0 1 1970
box -8 -3 16 105
use FILL  FILL_1314
timestamp 1714281807
transform 1 0 512 0 1 1970
box -8 -3 16 105
use FILL  FILL_1315
timestamp 1714281807
transform 1 0 472 0 1 1970
box -8 -3 16 105
use FILL  FILL_1316
timestamp 1714281807
transform 1 0 464 0 1 1970
box -8 -3 16 105
use FILL  FILL_1317
timestamp 1714281807
transform 1 0 456 0 1 1970
box -8 -3 16 105
use FILL  FILL_1318
timestamp 1714281807
transform 1 0 448 0 1 1970
box -8 -3 16 105
use FILL  FILL_1319
timestamp 1714281807
transform 1 0 440 0 1 1970
box -8 -3 16 105
use FILL  FILL_1320
timestamp 1714281807
transform 1 0 432 0 1 1970
box -8 -3 16 105
use FILL  FILL_1321
timestamp 1714281807
transform 1 0 424 0 1 1970
box -8 -3 16 105
use FILL  FILL_1322
timestamp 1714281807
transform 1 0 384 0 1 1970
box -8 -3 16 105
use FILL  FILL_1323
timestamp 1714281807
transform 1 0 376 0 1 1970
box -8 -3 16 105
use FILL  FILL_1324
timestamp 1714281807
transform 1 0 368 0 1 1970
box -8 -3 16 105
use FILL  FILL_1325
timestamp 1714281807
transform 1 0 360 0 1 1970
box -8 -3 16 105
use FILL  FILL_1326
timestamp 1714281807
transform 1 0 352 0 1 1970
box -8 -3 16 105
use FILL  FILL_1327
timestamp 1714281807
transform 1 0 344 0 1 1970
box -8 -3 16 105
use FILL  FILL_1328
timestamp 1714281807
transform 1 0 336 0 1 1970
box -8 -3 16 105
use FILL  FILL_1329
timestamp 1714281807
transform 1 0 328 0 1 1970
box -8 -3 16 105
use FILL  FILL_1330
timestamp 1714281807
transform 1 0 320 0 1 1970
box -8 -3 16 105
use FILL  FILL_1331
timestamp 1714281807
transform 1 0 296 0 1 1970
box -8 -3 16 105
use FILL  FILL_1332
timestamp 1714281807
transform 1 0 288 0 1 1970
box -8 -3 16 105
use FILL  FILL_1333
timestamp 1714281807
transform 1 0 280 0 1 1970
box -8 -3 16 105
use FILL  FILL_1334
timestamp 1714281807
transform 1 0 272 0 1 1970
box -8 -3 16 105
use FILL  FILL_1335
timestamp 1714281807
transform 1 0 264 0 1 1970
box -8 -3 16 105
use FILL  FILL_1336
timestamp 1714281807
transform 1 0 256 0 1 1970
box -8 -3 16 105
use FILL  FILL_1337
timestamp 1714281807
transform 1 0 248 0 1 1970
box -8 -3 16 105
use FILL  FILL_1338
timestamp 1714281807
transform 1 0 144 0 1 1970
box -8 -3 16 105
use FILL  FILL_1339
timestamp 1714281807
transform 1 0 136 0 1 1970
box -8 -3 16 105
use FILL  FILL_1340
timestamp 1714281807
transform 1 0 128 0 1 1970
box -8 -3 16 105
use FILL  FILL_1341
timestamp 1714281807
transform 1 0 120 0 1 1970
box -8 -3 16 105
use FILL  FILL_1342
timestamp 1714281807
transform 1 0 112 0 1 1970
box -8 -3 16 105
use FILL  FILL_1343
timestamp 1714281807
transform 1 0 104 0 1 1970
box -8 -3 16 105
use FILL  FILL_1344
timestamp 1714281807
transform 1 0 96 0 1 1970
box -8 -3 16 105
use FILL  FILL_1345
timestamp 1714281807
transform 1 0 88 0 1 1970
box -8 -3 16 105
use FILL  FILL_1346
timestamp 1714281807
transform 1 0 80 0 1 1970
box -8 -3 16 105
use FILL  FILL_1347
timestamp 1714281807
transform 1 0 72 0 1 1970
box -8 -3 16 105
use FILL  FILL_1348
timestamp 1714281807
transform 1 0 3000 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1349
timestamp 1714281807
transform 1 0 2992 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1350
timestamp 1714281807
transform 1 0 2984 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1351
timestamp 1714281807
transform 1 0 2976 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1352
timestamp 1714281807
transform 1 0 2968 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1353
timestamp 1714281807
transform 1 0 2864 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1354
timestamp 1714281807
transform 1 0 2856 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1355
timestamp 1714281807
transform 1 0 2848 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1356
timestamp 1714281807
transform 1 0 2816 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1357
timestamp 1714281807
transform 1 0 2808 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1358
timestamp 1714281807
transform 1 0 2784 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1359
timestamp 1714281807
transform 1 0 2776 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1360
timestamp 1714281807
transform 1 0 2768 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1361
timestamp 1714281807
transform 1 0 2760 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1362
timestamp 1714281807
transform 1 0 2720 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1363
timestamp 1714281807
transform 1 0 2712 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1364
timestamp 1714281807
transform 1 0 2608 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1365
timestamp 1714281807
transform 1 0 2600 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1366
timestamp 1714281807
transform 1 0 2592 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1367
timestamp 1714281807
transform 1 0 2584 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1368
timestamp 1714281807
transform 1 0 2576 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1369
timestamp 1714281807
transform 1 0 2528 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1370
timestamp 1714281807
transform 1 0 2520 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1371
timestamp 1714281807
transform 1 0 2416 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1372
timestamp 1714281807
transform 1 0 2408 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1373
timestamp 1714281807
transform 1 0 2400 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1374
timestamp 1714281807
transform 1 0 2360 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1375
timestamp 1714281807
transform 1 0 2296 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1376
timestamp 1714281807
transform 1 0 2288 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1377
timestamp 1714281807
transform 1 0 2280 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1378
timestamp 1714281807
transform 1 0 2272 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1379
timestamp 1714281807
transform 1 0 2224 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1380
timestamp 1714281807
transform 1 0 2216 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1381
timestamp 1714281807
transform 1 0 2208 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1382
timestamp 1714281807
transform 1 0 2104 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1383
timestamp 1714281807
transform 1 0 2080 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1384
timestamp 1714281807
transform 1 0 2072 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1385
timestamp 1714281807
transform 1 0 2064 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1386
timestamp 1714281807
transform 1 0 2056 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1387
timestamp 1714281807
transform 1 0 2024 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1388
timestamp 1714281807
transform 1 0 2016 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1389
timestamp 1714281807
transform 1 0 2008 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1390
timestamp 1714281807
transform 1 0 2000 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1391
timestamp 1714281807
transform 1 0 1992 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1392
timestamp 1714281807
transform 1 0 1984 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1393
timestamp 1714281807
transform 1 0 1952 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1394
timestamp 1714281807
transform 1 0 1944 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1395
timestamp 1714281807
transform 1 0 1936 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1396
timestamp 1714281807
transform 1 0 1928 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1397
timestamp 1714281807
transform 1 0 1920 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1398
timestamp 1714281807
transform 1 0 1912 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1399
timestamp 1714281807
transform 1 0 1904 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1400
timestamp 1714281807
transform 1 0 1872 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1401
timestamp 1714281807
transform 1 0 1808 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1402
timestamp 1714281807
transform 1 0 1704 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1403
timestamp 1714281807
transform 1 0 1600 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1404
timestamp 1714281807
transform 1 0 1568 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1405
timestamp 1714281807
transform 1 0 1560 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1406
timestamp 1714281807
transform 1 0 1552 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1407
timestamp 1714281807
transform 1 0 1448 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1408
timestamp 1714281807
transform 1 0 1424 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1409
timestamp 1714281807
transform 1 0 1416 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1410
timestamp 1714281807
transform 1 0 1408 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1411
timestamp 1714281807
transform 1 0 1400 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1412
timestamp 1714281807
transform 1 0 1352 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1413
timestamp 1714281807
transform 1 0 1344 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1414
timestamp 1714281807
transform 1 0 1336 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1415
timestamp 1714281807
transform 1 0 1328 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1416
timestamp 1714281807
transform 1 0 1320 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1417
timestamp 1714281807
transform 1 0 1312 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1418
timestamp 1714281807
transform 1 0 1264 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1419
timestamp 1714281807
transform 1 0 1256 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1420
timestamp 1714281807
transform 1 0 1248 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1421
timestamp 1714281807
transform 1 0 1224 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1422
timestamp 1714281807
transform 1 0 1216 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1423
timestamp 1714281807
transform 1 0 1208 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1424
timestamp 1714281807
transform 1 0 1184 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1425
timestamp 1714281807
transform 1 0 1176 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1426
timestamp 1714281807
transform 1 0 1168 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1427
timestamp 1714281807
transform 1 0 1128 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1428
timestamp 1714281807
transform 1 0 1120 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1429
timestamp 1714281807
transform 1 0 1112 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1430
timestamp 1714281807
transform 1 0 1104 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1431
timestamp 1714281807
transform 1 0 1096 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1432
timestamp 1714281807
transform 1 0 1072 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1433
timestamp 1714281807
transform 1 0 1064 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1434
timestamp 1714281807
transform 1 0 1032 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1435
timestamp 1714281807
transform 1 0 1024 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1436
timestamp 1714281807
transform 1 0 1016 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1437
timestamp 1714281807
transform 1 0 1008 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1438
timestamp 1714281807
transform 1 0 1000 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1439
timestamp 1714281807
transform 1 0 992 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1440
timestamp 1714281807
transform 1 0 960 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1441
timestamp 1714281807
transform 1 0 952 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1442
timestamp 1714281807
transform 1 0 944 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1443
timestamp 1714281807
transform 1 0 936 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1444
timestamp 1714281807
transform 1 0 928 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1445
timestamp 1714281807
transform 1 0 888 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1446
timestamp 1714281807
transform 1 0 880 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1447
timestamp 1714281807
transform 1 0 872 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1448
timestamp 1714281807
transform 1 0 864 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1449
timestamp 1714281807
transform 1 0 856 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1450
timestamp 1714281807
transform 1 0 848 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1451
timestamp 1714281807
transform 1 0 816 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1452
timestamp 1714281807
transform 1 0 808 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1453
timestamp 1714281807
transform 1 0 800 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1454
timestamp 1714281807
transform 1 0 792 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1455
timestamp 1714281807
transform 1 0 784 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1456
timestamp 1714281807
transform 1 0 776 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1457
timestamp 1714281807
transform 1 0 736 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1458
timestamp 1714281807
transform 1 0 728 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1459
timestamp 1714281807
transform 1 0 720 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1460
timestamp 1714281807
transform 1 0 712 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1461
timestamp 1714281807
transform 1 0 704 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1462
timestamp 1714281807
transform 1 0 696 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1463
timestamp 1714281807
transform 1 0 688 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1464
timestamp 1714281807
transform 1 0 680 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1465
timestamp 1714281807
transform 1 0 672 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1466
timestamp 1714281807
transform 1 0 624 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1467
timestamp 1714281807
transform 1 0 616 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1468
timestamp 1714281807
transform 1 0 608 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1469
timestamp 1714281807
transform 1 0 600 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1470
timestamp 1714281807
transform 1 0 592 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1471
timestamp 1714281807
transform 1 0 488 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1472
timestamp 1714281807
transform 1 0 480 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1473
timestamp 1714281807
transform 1 0 472 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1474
timestamp 1714281807
transform 1 0 368 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1475
timestamp 1714281807
transform 1 0 360 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1476
timestamp 1714281807
transform 1 0 352 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1477
timestamp 1714281807
transform 1 0 320 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1478
timestamp 1714281807
transform 1 0 312 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1479
timestamp 1714281807
transform 1 0 304 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1480
timestamp 1714281807
transform 1 0 296 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1481
timestamp 1714281807
transform 1 0 288 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1482
timestamp 1714281807
transform 1 0 280 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1483
timestamp 1714281807
transform 1 0 248 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1484
timestamp 1714281807
transform 1 0 240 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1485
timestamp 1714281807
transform 1 0 232 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1486
timestamp 1714281807
transform 1 0 224 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1487
timestamp 1714281807
transform 1 0 216 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1488
timestamp 1714281807
transform 1 0 192 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1489
timestamp 1714281807
transform 1 0 184 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1490
timestamp 1714281807
transform 1 0 176 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1491
timestamp 1714281807
transform 1 0 168 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1492
timestamp 1714281807
transform 1 0 160 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1493
timestamp 1714281807
transform 1 0 152 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1494
timestamp 1714281807
transform 1 0 144 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1495
timestamp 1714281807
transform 1 0 136 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1496
timestamp 1714281807
transform 1 0 128 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1497
timestamp 1714281807
transform 1 0 120 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1498
timestamp 1714281807
transform 1 0 112 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1499
timestamp 1714281807
transform 1 0 104 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1500
timestamp 1714281807
transform 1 0 96 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1501
timestamp 1714281807
transform 1 0 88 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1502
timestamp 1714281807
transform 1 0 80 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1503
timestamp 1714281807
transform 1 0 72 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1504
timestamp 1714281807
transform 1 0 3000 0 1 1770
box -8 -3 16 105
use FILL  FILL_1505
timestamp 1714281807
transform 1 0 2992 0 1 1770
box -8 -3 16 105
use FILL  FILL_1506
timestamp 1714281807
transform 1 0 2984 0 1 1770
box -8 -3 16 105
use FILL  FILL_1507
timestamp 1714281807
transform 1 0 2976 0 1 1770
box -8 -3 16 105
use FILL  FILL_1508
timestamp 1714281807
transform 1 0 2968 0 1 1770
box -8 -3 16 105
use FILL  FILL_1509
timestamp 1714281807
transform 1 0 2960 0 1 1770
box -8 -3 16 105
use FILL  FILL_1510
timestamp 1714281807
transform 1 0 2856 0 1 1770
box -8 -3 16 105
use FILL  FILL_1511
timestamp 1714281807
transform 1 0 2848 0 1 1770
box -8 -3 16 105
use FILL  FILL_1512
timestamp 1714281807
transform 1 0 2840 0 1 1770
box -8 -3 16 105
use FILL  FILL_1513
timestamp 1714281807
transform 1 0 2832 0 1 1770
box -8 -3 16 105
use FILL  FILL_1514
timestamp 1714281807
transform 1 0 2800 0 1 1770
box -8 -3 16 105
use FILL  FILL_1515
timestamp 1714281807
transform 1 0 2792 0 1 1770
box -8 -3 16 105
use FILL  FILL_1516
timestamp 1714281807
transform 1 0 2784 0 1 1770
box -8 -3 16 105
use FILL  FILL_1517
timestamp 1714281807
transform 1 0 2776 0 1 1770
box -8 -3 16 105
use FILL  FILL_1518
timestamp 1714281807
transform 1 0 2768 0 1 1770
box -8 -3 16 105
use FILL  FILL_1519
timestamp 1714281807
transform 1 0 2760 0 1 1770
box -8 -3 16 105
use FILL  FILL_1520
timestamp 1714281807
transform 1 0 2736 0 1 1770
box -8 -3 16 105
use FILL  FILL_1521
timestamp 1714281807
transform 1 0 2696 0 1 1770
box -8 -3 16 105
use FILL  FILL_1522
timestamp 1714281807
transform 1 0 2688 0 1 1770
box -8 -3 16 105
use FILL  FILL_1523
timestamp 1714281807
transform 1 0 2680 0 1 1770
box -8 -3 16 105
use FILL  FILL_1524
timestamp 1714281807
transform 1 0 2576 0 1 1770
box -8 -3 16 105
use FILL  FILL_1525
timestamp 1714281807
transform 1 0 2472 0 1 1770
box -8 -3 16 105
use FILL  FILL_1526
timestamp 1714281807
transform 1 0 2464 0 1 1770
box -8 -3 16 105
use FILL  FILL_1527
timestamp 1714281807
transform 1 0 2456 0 1 1770
box -8 -3 16 105
use FILL  FILL_1528
timestamp 1714281807
transform 1 0 2448 0 1 1770
box -8 -3 16 105
use FILL  FILL_1529
timestamp 1714281807
transform 1 0 2440 0 1 1770
box -8 -3 16 105
use FILL  FILL_1530
timestamp 1714281807
transform 1 0 2400 0 1 1770
box -8 -3 16 105
use FILL  FILL_1531
timestamp 1714281807
transform 1 0 2392 0 1 1770
box -8 -3 16 105
use FILL  FILL_1532
timestamp 1714281807
transform 1 0 2384 0 1 1770
box -8 -3 16 105
use FILL  FILL_1533
timestamp 1714281807
transform 1 0 2376 0 1 1770
box -8 -3 16 105
use FILL  FILL_1534
timestamp 1714281807
transform 1 0 2368 0 1 1770
box -8 -3 16 105
use FILL  FILL_1535
timestamp 1714281807
transform 1 0 2360 0 1 1770
box -8 -3 16 105
use FILL  FILL_1536
timestamp 1714281807
transform 1 0 2352 0 1 1770
box -8 -3 16 105
use FILL  FILL_1537
timestamp 1714281807
transform 1 0 2304 0 1 1770
box -8 -3 16 105
use FILL  FILL_1538
timestamp 1714281807
transform 1 0 2296 0 1 1770
box -8 -3 16 105
use FILL  FILL_1539
timestamp 1714281807
transform 1 0 2288 0 1 1770
box -8 -3 16 105
use FILL  FILL_1540
timestamp 1714281807
transform 1 0 2280 0 1 1770
box -8 -3 16 105
use FILL  FILL_1541
timestamp 1714281807
transform 1 0 2272 0 1 1770
box -8 -3 16 105
use FILL  FILL_1542
timestamp 1714281807
transform 1 0 2264 0 1 1770
box -8 -3 16 105
use FILL  FILL_1543
timestamp 1714281807
transform 1 0 2256 0 1 1770
box -8 -3 16 105
use FILL  FILL_1544
timestamp 1714281807
transform 1 0 2216 0 1 1770
box -8 -3 16 105
use FILL  FILL_1545
timestamp 1714281807
transform 1 0 2208 0 1 1770
box -8 -3 16 105
use FILL  FILL_1546
timestamp 1714281807
transform 1 0 2200 0 1 1770
box -8 -3 16 105
use FILL  FILL_1547
timestamp 1714281807
transform 1 0 2192 0 1 1770
box -8 -3 16 105
use FILL  FILL_1548
timestamp 1714281807
transform 1 0 2184 0 1 1770
box -8 -3 16 105
use FILL  FILL_1549
timestamp 1714281807
transform 1 0 2176 0 1 1770
box -8 -3 16 105
use FILL  FILL_1550
timestamp 1714281807
transform 1 0 2168 0 1 1770
box -8 -3 16 105
use FILL  FILL_1551
timestamp 1714281807
transform 1 0 2128 0 1 1770
box -8 -3 16 105
use FILL  FILL_1552
timestamp 1714281807
transform 1 0 2120 0 1 1770
box -8 -3 16 105
use FILL  FILL_1553
timestamp 1714281807
transform 1 0 2088 0 1 1770
box -8 -3 16 105
use FILL  FILL_1554
timestamp 1714281807
transform 1 0 2080 0 1 1770
box -8 -3 16 105
use FILL  FILL_1555
timestamp 1714281807
transform 1 0 1976 0 1 1770
box -8 -3 16 105
use FILL  FILL_1556
timestamp 1714281807
transform 1 0 1968 0 1 1770
box -8 -3 16 105
use FILL  FILL_1557
timestamp 1714281807
transform 1 0 1960 0 1 1770
box -8 -3 16 105
use FILL  FILL_1558
timestamp 1714281807
transform 1 0 1936 0 1 1770
box -8 -3 16 105
use FILL  FILL_1559
timestamp 1714281807
transform 1 0 1928 0 1 1770
box -8 -3 16 105
use FILL  FILL_1560
timestamp 1714281807
transform 1 0 1896 0 1 1770
box -8 -3 16 105
use FILL  FILL_1561
timestamp 1714281807
transform 1 0 1888 0 1 1770
box -8 -3 16 105
use FILL  FILL_1562
timestamp 1714281807
transform 1 0 1880 0 1 1770
box -8 -3 16 105
use FILL  FILL_1563
timestamp 1714281807
transform 1 0 1872 0 1 1770
box -8 -3 16 105
use FILL  FILL_1564
timestamp 1714281807
transform 1 0 1848 0 1 1770
box -8 -3 16 105
use FILL  FILL_1565
timestamp 1714281807
transform 1 0 1840 0 1 1770
box -8 -3 16 105
use FILL  FILL_1566
timestamp 1714281807
transform 1 0 1832 0 1 1770
box -8 -3 16 105
use FILL  FILL_1567
timestamp 1714281807
transform 1 0 1824 0 1 1770
box -8 -3 16 105
use FILL  FILL_1568
timestamp 1714281807
transform 1 0 1816 0 1 1770
box -8 -3 16 105
use FILL  FILL_1569
timestamp 1714281807
transform 1 0 1808 0 1 1770
box -8 -3 16 105
use FILL  FILL_1570
timestamp 1714281807
transform 1 0 1784 0 1 1770
box -8 -3 16 105
use FILL  FILL_1571
timestamp 1714281807
transform 1 0 1776 0 1 1770
box -8 -3 16 105
use FILL  FILL_1572
timestamp 1714281807
transform 1 0 1768 0 1 1770
box -8 -3 16 105
use FILL  FILL_1573
timestamp 1714281807
transform 1 0 1760 0 1 1770
box -8 -3 16 105
use FILL  FILL_1574
timestamp 1714281807
transform 1 0 1728 0 1 1770
box -8 -3 16 105
use FILL  FILL_1575
timestamp 1714281807
transform 1 0 1720 0 1 1770
box -8 -3 16 105
use FILL  FILL_1576
timestamp 1714281807
transform 1 0 1712 0 1 1770
box -8 -3 16 105
use FILL  FILL_1577
timestamp 1714281807
transform 1 0 1704 0 1 1770
box -8 -3 16 105
use FILL  FILL_1578
timestamp 1714281807
transform 1 0 1696 0 1 1770
box -8 -3 16 105
use FILL  FILL_1579
timestamp 1714281807
transform 1 0 1688 0 1 1770
box -8 -3 16 105
use FILL  FILL_1580
timestamp 1714281807
transform 1 0 1680 0 1 1770
box -8 -3 16 105
use FILL  FILL_1581
timestamp 1714281807
transform 1 0 1672 0 1 1770
box -8 -3 16 105
use FILL  FILL_1582
timestamp 1714281807
transform 1 0 1664 0 1 1770
box -8 -3 16 105
use FILL  FILL_1583
timestamp 1714281807
transform 1 0 1656 0 1 1770
box -8 -3 16 105
use FILL  FILL_1584
timestamp 1714281807
transform 1 0 1648 0 1 1770
box -8 -3 16 105
use FILL  FILL_1585
timestamp 1714281807
transform 1 0 1640 0 1 1770
box -8 -3 16 105
use FILL  FILL_1586
timestamp 1714281807
transform 1 0 1616 0 1 1770
box -8 -3 16 105
use FILL  FILL_1587
timestamp 1714281807
transform 1 0 1608 0 1 1770
box -8 -3 16 105
use FILL  FILL_1588
timestamp 1714281807
transform 1 0 1504 0 1 1770
box -8 -3 16 105
use FILL  FILL_1589
timestamp 1714281807
transform 1 0 1496 0 1 1770
box -8 -3 16 105
use FILL  FILL_1590
timestamp 1714281807
transform 1 0 1488 0 1 1770
box -8 -3 16 105
use FILL  FILL_1591
timestamp 1714281807
transform 1 0 1480 0 1 1770
box -8 -3 16 105
use FILL  FILL_1592
timestamp 1714281807
transform 1 0 1376 0 1 1770
box -8 -3 16 105
use FILL  FILL_1593
timestamp 1714281807
transform 1 0 1368 0 1 1770
box -8 -3 16 105
use FILL  FILL_1594
timestamp 1714281807
transform 1 0 1360 0 1 1770
box -8 -3 16 105
use FILL  FILL_1595
timestamp 1714281807
transform 1 0 1336 0 1 1770
box -8 -3 16 105
use FILL  FILL_1596
timestamp 1714281807
transform 1 0 1328 0 1 1770
box -8 -3 16 105
use FILL  FILL_1597
timestamp 1714281807
transform 1 0 1320 0 1 1770
box -8 -3 16 105
use FILL  FILL_1598
timestamp 1714281807
transform 1 0 1312 0 1 1770
box -8 -3 16 105
use FILL  FILL_1599
timestamp 1714281807
transform 1 0 1272 0 1 1770
box -8 -3 16 105
use FILL  FILL_1600
timestamp 1714281807
transform 1 0 1264 0 1 1770
box -8 -3 16 105
use FILL  FILL_1601
timestamp 1714281807
transform 1 0 1256 0 1 1770
box -8 -3 16 105
use FILL  FILL_1602
timestamp 1714281807
transform 1 0 1248 0 1 1770
box -8 -3 16 105
use FILL  FILL_1603
timestamp 1714281807
transform 1 0 1240 0 1 1770
box -8 -3 16 105
use FILL  FILL_1604
timestamp 1714281807
transform 1 0 1232 0 1 1770
box -8 -3 16 105
use FILL  FILL_1605
timestamp 1714281807
transform 1 0 1200 0 1 1770
box -8 -3 16 105
use FILL  FILL_1606
timestamp 1714281807
transform 1 0 1192 0 1 1770
box -8 -3 16 105
use FILL  FILL_1607
timestamp 1714281807
transform 1 0 1184 0 1 1770
box -8 -3 16 105
use FILL  FILL_1608
timestamp 1714281807
transform 1 0 1080 0 1 1770
box -8 -3 16 105
use FILL  FILL_1609
timestamp 1714281807
transform 1 0 1072 0 1 1770
box -8 -3 16 105
use FILL  FILL_1610
timestamp 1714281807
transform 1 0 1064 0 1 1770
box -8 -3 16 105
use FILL  FILL_1611
timestamp 1714281807
transform 1 0 1056 0 1 1770
box -8 -3 16 105
use FILL  FILL_1612
timestamp 1714281807
transform 1 0 1048 0 1 1770
box -8 -3 16 105
use FILL  FILL_1613
timestamp 1714281807
transform 1 0 1040 0 1 1770
box -8 -3 16 105
use FILL  FILL_1614
timestamp 1714281807
transform 1 0 984 0 1 1770
box -8 -3 16 105
use FILL  FILL_1615
timestamp 1714281807
transform 1 0 976 0 1 1770
box -8 -3 16 105
use FILL  FILL_1616
timestamp 1714281807
transform 1 0 968 0 1 1770
box -8 -3 16 105
use FILL  FILL_1617
timestamp 1714281807
transform 1 0 960 0 1 1770
box -8 -3 16 105
use FILL  FILL_1618
timestamp 1714281807
transform 1 0 952 0 1 1770
box -8 -3 16 105
use FILL  FILL_1619
timestamp 1714281807
transform 1 0 928 0 1 1770
box -8 -3 16 105
use FILL  FILL_1620
timestamp 1714281807
transform 1 0 920 0 1 1770
box -8 -3 16 105
use FILL  FILL_1621
timestamp 1714281807
transform 1 0 912 0 1 1770
box -8 -3 16 105
use FILL  FILL_1622
timestamp 1714281807
transform 1 0 904 0 1 1770
box -8 -3 16 105
use FILL  FILL_1623
timestamp 1714281807
transform 1 0 896 0 1 1770
box -8 -3 16 105
use FILL  FILL_1624
timestamp 1714281807
transform 1 0 888 0 1 1770
box -8 -3 16 105
use FILL  FILL_1625
timestamp 1714281807
transform 1 0 840 0 1 1770
box -8 -3 16 105
use FILL  FILL_1626
timestamp 1714281807
transform 1 0 832 0 1 1770
box -8 -3 16 105
use FILL  FILL_1627
timestamp 1714281807
transform 1 0 824 0 1 1770
box -8 -3 16 105
use FILL  FILL_1628
timestamp 1714281807
transform 1 0 816 0 1 1770
box -8 -3 16 105
use FILL  FILL_1629
timestamp 1714281807
transform 1 0 808 0 1 1770
box -8 -3 16 105
use FILL  FILL_1630
timestamp 1714281807
transform 1 0 800 0 1 1770
box -8 -3 16 105
use FILL  FILL_1631
timestamp 1714281807
transform 1 0 792 0 1 1770
box -8 -3 16 105
use FILL  FILL_1632
timestamp 1714281807
transform 1 0 768 0 1 1770
box -8 -3 16 105
use FILL  FILL_1633
timestamp 1714281807
transform 1 0 760 0 1 1770
box -8 -3 16 105
use FILL  FILL_1634
timestamp 1714281807
transform 1 0 752 0 1 1770
box -8 -3 16 105
use FILL  FILL_1635
timestamp 1714281807
transform 1 0 720 0 1 1770
box -8 -3 16 105
use FILL  FILL_1636
timestamp 1714281807
transform 1 0 712 0 1 1770
box -8 -3 16 105
use FILL  FILL_1637
timestamp 1714281807
transform 1 0 704 0 1 1770
box -8 -3 16 105
use FILL  FILL_1638
timestamp 1714281807
transform 1 0 696 0 1 1770
box -8 -3 16 105
use FILL  FILL_1639
timestamp 1714281807
transform 1 0 688 0 1 1770
box -8 -3 16 105
use FILL  FILL_1640
timestamp 1714281807
transform 1 0 680 0 1 1770
box -8 -3 16 105
use FILL  FILL_1641
timestamp 1714281807
transform 1 0 640 0 1 1770
box -8 -3 16 105
use FILL  FILL_1642
timestamp 1714281807
transform 1 0 632 0 1 1770
box -8 -3 16 105
use FILL  FILL_1643
timestamp 1714281807
transform 1 0 608 0 1 1770
box -8 -3 16 105
use FILL  FILL_1644
timestamp 1714281807
transform 1 0 600 0 1 1770
box -8 -3 16 105
use FILL  FILL_1645
timestamp 1714281807
transform 1 0 592 0 1 1770
box -8 -3 16 105
use FILL  FILL_1646
timestamp 1714281807
transform 1 0 584 0 1 1770
box -8 -3 16 105
use FILL  FILL_1647
timestamp 1714281807
transform 1 0 576 0 1 1770
box -8 -3 16 105
use FILL  FILL_1648
timestamp 1714281807
transform 1 0 536 0 1 1770
box -8 -3 16 105
use FILL  FILL_1649
timestamp 1714281807
transform 1 0 528 0 1 1770
box -8 -3 16 105
use FILL  FILL_1650
timestamp 1714281807
transform 1 0 520 0 1 1770
box -8 -3 16 105
use FILL  FILL_1651
timestamp 1714281807
transform 1 0 488 0 1 1770
box -8 -3 16 105
use FILL  FILL_1652
timestamp 1714281807
transform 1 0 480 0 1 1770
box -8 -3 16 105
use FILL  FILL_1653
timestamp 1714281807
transform 1 0 472 0 1 1770
box -8 -3 16 105
use FILL  FILL_1654
timestamp 1714281807
transform 1 0 464 0 1 1770
box -8 -3 16 105
use FILL  FILL_1655
timestamp 1714281807
transform 1 0 456 0 1 1770
box -8 -3 16 105
use FILL  FILL_1656
timestamp 1714281807
transform 1 0 448 0 1 1770
box -8 -3 16 105
use FILL  FILL_1657
timestamp 1714281807
transform 1 0 400 0 1 1770
box -8 -3 16 105
use FILL  FILL_1658
timestamp 1714281807
transform 1 0 392 0 1 1770
box -8 -3 16 105
use FILL  FILL_1659
timestamp 1714281807
transform 1 0 384 0 1 1770
box -8 -3 16 105
use FILL  FILL_1660
timestamp 1714281807
transform 1 0 280 0 1 1770
box -8 -3 16 105
use FILL  FILL_1661
timestamp 1714281807
transform 1 0 272 0 1 1770
box -8 -3 16 105
use FILL  FILL_1662
timestamp 1714281807
transform 1 0 232 0 1 1770
box -8 -3 16 105
use FILL  FILL_1663
timestamp 1714281807
transform 1 0 224 0 1 1770
box -8 -3 16 105
use FILL  FILL_1664
timestamp 1714281807
transform 1 0 216 0 1 1770
box -8 -3 16 105
use FILL  FILL_1665
timestamp 1714281807
transform 1 0 208 0 1 1770
box -8 -3 16 105
use FILL  FILL_1666
timestamp 1714281807
transform 1 0 184 0 1 1770
box -8 -3 16 105
use FILL  FILL_1667
timestamp 1714281807
transform 1 0 80 0 1 1770
box -8 -3 16 105
use FILL  FILL_1668
timestamp 1714281807
transform 1 0 72 0 1 1770
box -8 -3 16 105
use FILL  FILL_1669
timestamp 1714281807
transform 1 0 3000 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1670
timestamp 1714281807
transform 1 0 2992 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1671
timestamp 1714281807
transform 1 0 2984 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1672
timestamp 1714281807
transform 1 0 2976 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1673
timestamp 1714281807
transform 1 0 2968 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1674
timestamp 1714281807
transform 1 0 2960 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1675
timestamp 1714281807
transform 1 0 2856 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1676
timestamp 1714281807
transform 1 0 2848 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1677
timestamp 1714281807
transform 1 0 2840 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1678
timestamp 1714281807
transform 1 0 2808 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1679
timestamp 1714281807
transform 1 0 2800 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1680
timestamp 1714281807
transform 1 0 2792 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1681
timestamp 1714281807
transform 1 0 2784 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1682
timestamp 1714281807
transform 1 0 2760 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1683
timestamp 1714281807
transform 1 0 2752 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1684
timestamp 1714281807
transform 1 0 2712 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1685
timestamp 1714281807
transform 1 0 2704 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1686
timestamp 1714281807
transform 1 0 2696 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1687
timestamp 1714281807
transform 1 0 2592 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1688
timestamp 1714281807
transform 1 0 2488 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1689
timestamp 1714281807
transform 1 0 2480 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1690
timestamp 1714281807
transform 1 0 2448 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1691
timestamp 1714281807
transform 1 0 2440 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1692
timestamp 1714281807
transform 1 0 2432 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1693
timestamp 1714281807
transform 1 0 2328 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1694
timestamp 1714281807
transform 1 0 2320 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1695
timestamp 1714281807
transform 1 0 2312 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1696
timestamp 1714281807
transform 1 0 2232 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1697
timestamp 1714281807
transform 1 0 2224 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1698
timestamp 1714281807
transform 1 0 2216 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1699
timestamp 1714281807
transform 1 0 2208 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1700
timestamp 1714281807
transform 1 0 2200 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1701
timestamp 1714281807
transform 1 0 2192 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1702
timestamp 1714281807
transform 1 0 2184 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1703
timestamp 1714281807
transform 1 0 2176 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1704
timestamp 1714281807
transform 1 0 2168 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1705
timestamp 1714281807
transform 1 0 2128 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1706
timestamp 1714281807
transform 1 0 2120 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1707
timestamp 1714281807
transform 1 0 2112 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1708
timestamp 1714281807
transform 1 0 2008 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1709
timestamp 1714281807
transform 1 0 2000 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1710
timestamp 1714281807
transform 1 0 1896 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1711
timestamp 1714281807
transform 1 0 1792 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1712
timestamp 1714281807
transform 1 0 1784 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1713
timestamp 1714281807
transform 1 0 1776 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1714
timestamp 1714281807
transform 1 0 1768 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1715
timestamp 1714281807
transform 1 0 1728 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1716
timestamp 1714281807
transform 1 0 1720 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1717
timestamp 1714281807
transform 1 0 1712 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1718
timestamp 1714281807
transform 1 0 1704 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1719
timestamp 1714281807
transform 1 0 1696 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1720
timestamp 1714281807
transform 1 0 1688 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1721
timestamp 1714281807
transform 1 0 1680 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1722
timestamp 1714281807
transform 1 0 1632 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1723
timestamp 1714281807
transform 1 0 1624 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1724
timestamp 1714281807
transform 1 0 1616 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1725
timestamp 1714281807
transform 1 0 1608 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1726
timestamp 1714281807
transform 1 0 1600 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1727
timestamp 1714281807
transform 1 0 1592 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1728
timestamp 1714281807
transform 1 0 1584 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1729
timestamp 1714281807
transform 1 0 1544 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1730
timestamp 1714281807
transform 1 0 1536 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1731
timestamp 1714281807
transform 1 0 1528 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1732
timestamp 1714281807
transform 1 0 1520 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1733
timestamp 1714281807
transform 1 0 1512 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1734
timestamp 1714281807
transform 1 0 1408 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1735
timestamp 1714281807
transform 1 0 1400 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1736
timestamp 1714281807
transform 1 0 1392 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1737
timestamp 1714281807
transform 1 0 1288 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1738
timestamp 1714281807
transform 1 0 1280 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1739
timestamp 1714281807
transform 1 0 1272 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1740
timestamp 1714281807
transform 1 0 1240 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1741
timestamp 1714281807
transform 1 0 1232 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1742
timestamp 1714281807
transform 1 0 1224 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1743
timestamp 1714281807
transform 1 0 1216 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1744
timestamp 1714281807
transform 1 0 1208 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1745
timestamp 1714281807
transform 1 0 1184 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1746
timestamp 1714281807
transform 1 0 1160 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1747
timestamp 1714281807
transform 1 0 1152 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1748
timestamp 1714281807
transform 1 0 1144 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1749
timestamp 1714281807
transform 1 0 1136 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1750
timestamp 1714281807
transform 1 0 1128 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1751
timestamp 1714281807
transform 1 0 1080 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1752
timestamp 1714281807
transform 1 0 1072 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1753
timestamp 1714281807
transform 1 0 1064 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1754
timestamp 1714281807
transform 1 0 1056 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1755
timestamp 1714281807
transform 1 0 1048 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1756
timestamp 1714281807
transform 1 0 1024 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1757
timestamp 1714281807
transform 1 0 1016 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1758
timestamp 1714281807
transform 1 0 976 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1759
timestamp 1714281807
transform 1 0 968 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1760
timestamp 1714281807
transform 1 0 928 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1761
timestamp 1714281807
transform 1 0 920 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1762
timestamp 1714281807
transform 1 0 912 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1763
timestamp 1714281807
transform 1 0 904 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1764
timestamp 1714281807
transform 1 0 896 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1765
timestamp 1714281807
transform 1 0 848 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1766
timestamp 1714281807
transform 1 0 840 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1767
timestamp 1714281807
transform 1 0 832 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1768
timestamp 1714281807
transform 1 0 824 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1769
timestamp 1714281807
transform 1 0 816 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1770
timestamp 1714281807
transform 1 0 696 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1771
timestamp 1714281807
transform 1 0 688 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1772
timestamp 1714281807
transform 1 0 680 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1773
timestamp 1714281807
transform 1 0 672 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1774
timestamp 1714281807
transform 1 0 616 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1775
timestamp 1714281807
transform 1 0 608 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1776
timestamp 1714281807
transform 1 0 600 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1777
timestamp 1714281807
transform 1 0 592 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1778
timestamp 1714281807
transform 1 0 584 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1779
timestamp 1714281807
transform 1 0 576 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1780
timestamp 1714281807
transform 1 0 568 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1781
timestamp 1714281807
transform 1 0 560 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1782
timestamp 1714281807
transform 1 0 520 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1783
timestamp 1714281807
transform 1 0 512 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1784
timestamp 1714281807
transform 1 0 504 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1785
timestamp 1714281807
transform 1 0 496 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1786
timestamp 1714281807
transform 1 0 488 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1787
timestamp 1714281807
transform 1 0 464 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1788
timestamp 1714281807
transform 1 0 456 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1789
timestamp 1714281807
transform 1 0 448 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1790
timestamp 1714281807
transform 1 0 440 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1791
timestamp 1714281807
transform 1 0 432 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1792
timestamp 1714281807
transform 1 0 424 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1793
timestamp 1714281807
transform 1 0 384 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1794
timestamp 1714281807
transform 1 0 376 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1795
timestamp 1714281807
transform 1 0 368 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1796
timestamp 1714281807
transform 1 0 360 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1797
timestamp 1714281807
transform 1 0 256 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1798
timestamp 1714281807
transform 1 0 248 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1799
timestamp 1714281807
transform 1 0 240 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1800
timestamp 1714281807
transform 1 0 232 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1801
timestamp 1714281807
transform 1 0 224 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1802
timestamp 1714281807
transform 1 0 216 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1803
timestamp 1714281807
transform 1 0 208 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1804
timestamp 1714281807
transform 1 0 200 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1805
timestamp 1714281807
transform 1 0 192 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1806
timestamp 1714281807
transform 1 0 184 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1807
timestamp 1714281807
transform 1 0 176 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1808
timestamp 1714281807
transform 1 0 168 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1809
timestamp 1714281807
transform 1 0 160 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1810
timestamp 1714281807
transform 1 0 152 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1811
timestamp 1714281807
transform 1 0 144 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1812
timestamp 1714281807
transform 1 0 136 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1813
timestamp 1714281807
transform 1 0 128 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1814
timestamp 1714281807
transform 1 0 120 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1815
timestamp 1714281807
transform 1 0 112 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1816
timestamp 1714281807
transform 1 0 104 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1817
timestamp 1714281807
transform 1 0 96 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1818
timestamp 1714281807
transform 1 0 88 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1819
timestamp 1714281807
transform 1 0 80 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1820
timestamp 1714281807
transform 1 0 72 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1821
timestamp 1714281807
transform 1 0 3000 0 1 1570
box -8 -3 16 105
use FILL  FILL_1822
timestamp 1714281807
transform 1 0 2992 0 1 1570
box -8 -3 16 105
use FILL  FILL_1823
timestamp 1714281807
transform 1 0 2984 0 1 1570
box -8 -3 16 105
use FILL  FILL_1824
timestamp 1714281807
transform 1 0 2976 0 1 1570
box -8 -3 16 105
use FILL  FILL_1825
timestamp 1714281807
transform 1 0 2968 0 1 1570
box -8 -3 16 105
use FILL  FILL_1826
timestamp 1714281807
transform 1 0 2864 0 1 1570
box -8 -3 16 105
use FILL  FILL_1827
timestamp 1714281807
transform 1 0 2856 0 1 1570
box -8 -3 16 105
use FILL  FILL_1828
timestamp 1714281807
transform 1 0 2848 0 1 1570
box -8 -3 16 105
use FILL  FILL_1829
timestamp 1714281807
transform 1 0 2840 0 1 1570
box -8 -3 16 105
use FILL  FILL_1830
timestamp 1714281807
transform 1 0 2792 0 1 1570
box -8 -3 16 105
use FILL  FILL_1831
timestamp 1714281807
transform 1 0 2784 0 1 1570
box -8 -3 16 105
use FILL  FILL_1832
timestamp 1714281807
transform 1 0 2776 0 1 1570
box -8 -3 16 105
use FILL  FILL_1833
timestamp 1714281807
transform 1 0 2672 0 1 1570
box -8 -3 16 105
use FILL  FILL_1834
timestamp 1714281807
transform 1 0 2632 0 1 1570
box -8 -3 16 105
use FILL  FILL_1835
timestamp 1714281807
transform 1 0 2624 0 1 1570
box -8 -3 16 105
use FILL  FILL_1836
timestamp 1714281807
transform 1 0 2496 0 1 1570
box -8 -3 16 105
use FILL  FILL_1837
timestamp 1714281807
transform 1 0 2488 0 1 1570
box -8 -3 16 105
use FILL  FILL_1838
timestamp 1714281807
transform 1 0 2384 0 1 1570
box -8 -3 16 105
use FILL  FILL_1839
timestamp 1714281807
transform 1 0 2376 0 1 1570
box -8 -3 16 105
use FILL  FILL_1840
timestamp 1714281807
transform 1 0 2336 0 1 1570
box -8 -3 16 105
use FILL  FILL_1841
timestamp 1714281807
transform 1 0 2328 0 1 1570
box -8 -3 16 105
use FILL  FILL_1842
timestamp 1714281807
transform 1 0 2320 0 1 1570
box -8 -3 16 105
use FILL  FILL_1843
timestamp 1714281807
transform 1 0 2312 0 1 1570
box -8 -3 16 105
use FILL  FILL_1844
timestamp 1714281807
transform 1 0 2304 0 1 1570
box -8 -3 16 105
use FILL  FILL_1845
timestamp 1714281807
transform 1 0 2256 0 1 1570
box -8 -3 16 105
use FILL  FILL_1846
timestamp 1714281807
transform 1 0 2248 0 1 1570
box -8 -3 16 105
use FILL  FILL_1847
timestamp 1714281807
transform 1 0 2240 0 1 1570
box -8 -3 16 105
use FILL  FILL_1848
timestamp 1714281807
transform 1 0 2136 0 1 1570
box -8 -3 16 105
use FILL  FILL_1849
timestamp 1714281807
transform 1 0 2128 0 1 1570
box -8 -3 16 105
use FILL  FILL_1850
timestamp 1714281807
transform 1 0 2120 0 1 1570
box -8 -3 16 105
use FILL  FILL_1851
timestamp 1714281807
transform 1 0 2112 0 1 1570
box -8 -3 16 105
use FILL  FILL_1852
timestamp 1714281807
transform 1 0 2080 0 1 1570
box -8 -3 16 105
use FILL  FILL_1853
timestamp 1714281807
transform 1 0 2072 0 1 1570
box -8 -3 16 105
use FILL  FILL_1854
timestamp 1714281807
transform 1 0 2048 0 1 1570
box -8 -3 16 105
use FILL  FILL_1855
timestamp 1714281807
transform 1 0 2040 0 1 1570
box -8 -3 16 105
use FILL  FILL_1856
timestamp 1714281807
transform 1 0 2032 0 1 1570
box -8 -3 16 105
use FILL  FILL_1857
timestamp 1714281807
transform 1 0 2024 0 1 1570
box -8 -3 16 105
use FILL  FILL_1858
timestamp 1714281807
transform 1 0 2016 0 1 1570
box -8 -3 16 105
use FILL  FILL_1859
timestamp 1714281807
transform 1 0 2008 0 1 1570
box -8 -3 16 105
use FILL  FILL_1860
timestamp 1714281807
transform 1 0 1968 0 1 1570
box -8 -3 16 105
use FILL  FILL_1861
timestamp 1714281807
transform 1 0 1960 0 1 1570
box -8 -3 16 105
use FILL  FILL_1862
timestamp 1714281807
transform 1 0 1952 0 1 1570
box -8 -3 16 105
use FILL  FILL_1863
timestamp 1714281807
transform 1 0 1928 0 1 1570
box -8 -3 16 105
use FILL  FILL_1864
timestamp 1714281807
transform 1 0 1920 0 1 1570
box -8 -3 16 105
use FILL  FILL_1865
timestamp 1714281807
transform 1 0 1912 0 1 1570
box -8 -3 16 105
use FILL  FILL_1866
timestamp 1714281807
transform 1 0 1904 0 1 1570
box -8 -3 16 105
use FILL  FILL_1867
timestamp 1714281807
transform 1 0 1872 0 1 1570
box -8 -3 16 105
use FILL  FILL_1868
timestamp 1714281807
transform 1 0 1864 0 1 1570
box -8 -3 16 105
use FILL  FILL_1869
timestamp 1714281807
transform 1 0 1856 0 1 1570
box -8 -3 16 105
use FILL  FILL_1870
timestamp 1714281807
transform 1 0 1792 0 1 1570
box -8 -3 16 105
use FILL  FILL_1871
timestamp 1714281807
transform 1 0 1784 0 1 1570
box -8 -3 16 105
use FILL  FILL_1872
timestamp 1714281807
transform 1 0 1776 0 1 1570
box -8 -3 16 105
use FILL  FILL_1873
timestamp 1714281807
transform 1 0 1768 0 1 1570
box -8 -3 16 105
use FILL  FILL_1874
timestamp 1714281807
transform 1 0 1720 0 1 1570
box -8 -3 16 105
use FILL  FILL_1875
timestamp 1714281807
transform 1 0 1712 0 1 1570
box -8 -3 16 105
use FILL  FILL_1876
timestamp 1714281807
transform 1 0 1704 0 1 1570
box -8 -3 16 105
use FILL  FILL_1877
timestamp 1714281807
transform 1 0 1664 0 1 1570
box -8 -3 16 105
use FILL  FILL_1878
timestamp 1714281807
transform 1 0 1504 0 1 1570
box -8 -3 16 105
use FILL  FILL_1879
timestamp 1714281807
transform 1 0 1496 0 1 1570
box -8 -3 16 105
use FILL  FILL_1880
timestamp 1714281807
transform 1 0 1464 0 1 1570
box -8 -3 16 105
use FILL  FILL_1881
timestamp 1714281807
transform 1 0 1456 0 1 1570
box -8 -3 16 105
use FILL  FILL_1882
timestamp 1714281807
transform 1 0 1432 0 1 1570
box -8 -3 16 105
use FILL  FILL_1883
timestamp 1714281807
transform 1 0 1424 0 1 1570
box -8 -3 16 105
use FILL  FILL_1884
timestamp 1714281807
transform 1 0 1392 0 1 1570
box -8 -3 16 105
use FILL  FILL_1885
timestamp 1714281807
transform 1 0 1384 0 1 1570
box -8 -3 16 105
use FILL  FILL_1886
timestamp 1714281807
transform 1 0 1248 0 1 1570
box -8 -3 16 105
use FILL  FILL_1887
timestamp 1714281807
transform 1 0 1240 0 1 1570
box -8 -3 16 105
use FILL  FILL_1888
timestamp 1714281807
transform 1 0 1232 0 1 1570
box -8 -3 16 105
use FILL  FILL_1889
timestamp 1714281807
transform 1 0 1224 0 1 1570
box -8 -3 16 105
use FILL  FILL_1890
timestamp 1714281807
transform 1 0 1176 0 1 1570
box -8 -3 16 105
use FILL  FILL_1891
timestamp 1714281807
transform 1 0 1168 0 1 1570
box -8 -3 16 105
use FILL  FILL_1892
timestamp 1714281807
transform 1 0 1160 0 1 1570
box -8 -3 16 105
use FILL  FILL_1893
timestamp 1714281807
transform 1 0 1152 0 1 1570
box -8 -3 16 105
use FILL  FILL_1894
timestamp 1714281807
transform 1 0 1144 0 1 1570
box -8 -3 16 105
use FILL  FILL_1895
timestamp 1714281807
transform 1 0 1136 0 1 1570
box -8 -3 16 105
use FILL  FILL_1896
timestamp 1714281807
transform 1 0 1088 0 1 1570
box -8 -3 16 105
use FILL  FILL_1897
timestamp 1714281807
transform 1 0 1064 0 1 1570
box -8 -3 16 105
use FILL  FILL_1898
timestamp 1714281807
transform 1 0 1056 0 1 1570
box -8 -3 16 105
use FILL  FILL_1899
timestamp 1714281807
transform 1 0 1048 0 1 1570
box -8 -3 16 105
use FILL  FILL_1900
timestamp 1714281807
transform 1 0 1040 0 1 1570
box -8 -3 16 105
use FILL  FILL_1901
timestamp 1714281807
transform 1 0 1032 0 1 1570
box -8 -3 16 105
use FILL  FILL_1902
timestamp 1714281807
transform 1 0 984 0 1 1570
box -8 -3 16 105
use FILL  FILL_1903
timestamp 1714281807
transform 1 0 976 0 1 1570
box -8 -3 16 105
use FILL  FILL_1904
timestamp 1714281807
transform 1 0 968 0 1 1570
box -8 -3 16 105
use FILL  FILL_1905
timestamp 1714281807
transform 1 0 960 0 1 1570
box -8 -3 16 105
use FILL  FILL_1906
timestamp 1714281807
transform 1 0 952 0 1 1570
box -8 -3 16 105
use FILL  FILL_1907
timestamp 1714281807
transform 1 0 912 0 1 1570
box -8 -3 16 105
use FILL  FILL_1908
timestamp 1714281807
transform 1 0 904 0 1 1570
box -8 -3 16 105
use FILL  FILL_1909
timestamp 1714281807
transform 1 0 896 0 1 1570
box -8 -3 16 105
use FILL  FILL_1910
timestamp 1714281807
transform 1 0 888 0 1 1570
box -8 -3 16 105
use FILL  FILL_1911
timestamp 1714281807
transform 1 0 848 0 1 1570
box -8 -3 16 105
use FILL  FILL_1912
timestamp 1714281807
transform 1 0 840 0 1 1570
box -8 -3 16 105
use FILL  FILL_1913
timestamp 1714281807
transform 1 0 832 0 1 1570
box -8 -3 16 105
use FILL  FILL_1914
timestamp 1714281807
transform 1 0 800 0 1 1570
box -8 -3 16 105
use FILL  FILL_1915
timestamp 1714281807
transform 1 0 792 0 1 1570
box -8 -3 16 105
use FILL  FILL_1916
timestamp 1714281807
transform 1 0 784 0 1 1570
box -8 -3 16 105
use FILL  FILL_1917
timestamp 1714281807
transform 1 0 776 0 1 1570
box -8 -3 16 105
use FILL  FILL_1918
timestamp 1714281807
transform 1 0 768 0 1 1570
box -8 -3 16 105
use FILL  FILL_1919
timestamp 1714281807
transform 1 0 744 0 1 1570
box -8 -3 16 105
use FILL  FILL_1920
timestamp 1714281807
transform 1 0 704 0 1 1570
box -8 -3 16 105
use FILL  FILL_1921
timestamp 1714281807
transform 1 0 696 0 1 1570
box -8 -3 16 105
use FILL  FILL_1922
timestamp 1714281807
transform 1 0 688 0 1 1570
box -8 -3 16 105
use FILL  FILL_1923
timestamp 1714281807
transform 1 0 680 0 1 1570
box -8 -3 16 105
use FILL  FILL_1924
timestamp 1714281807
transform 1 0 672 0 1 1570
box -8 -3 16 105
use FILL  FILL_1925
timestamp 1714281807
transform 1 0 632 0 1 1570
box -8 -3 16 105
use FILL  FILL_1926
timestamp 1714281807
transform 1 0 624 0 1 1570
box -8 -3 16 105
use FILL  FILL_1927
timestamp 1714281807
transform 1 0 616 0 1 1570
box -8 -3 16 105
use FILL  FILL_1928
timestamp 1714281807
transform 1 0 608 0 1 1570
box -8 -3 16 105
use FILL  FILL_1929
timestamp 1714281807
transform 1 0 568 0 1 1570
box -8 -3 16 105
use FILL  FILL_1930
timestamp 1714281807
transform 1 0 560 0 1 1570
box -8 -3 16 105
use FILL  FILL_1931
timestamp 1714281807
transform 1 0 552 0 1 1570
box -8 -3 16 105
use FILL  FILL_1932
timestamp 1714281807
transform 1 0 544 0 1 1570
box -8 -3 16 105
use FILL  FILL_1933
timestamp 1714281807
transform 1 0 536 0 1 1570
box -8 -3 16 105
use FILL  FILL_1934
timestamp 1714281807
transform 1 0 496 0 1 1570
box -8 -3 16 105
use FILL  FILL_1935
timestamp 1714281807
transform 1 0 488 0 1 1570
box -8 -3 16 105
use FILL  FILL_1936
timestamp 1714281807
transform 1 0 480 0 1 1570
box -8 -3 16 105
use FILL  FILL_1937
timestamp 1714281807
transform 1 0 472 0 1 1570
box -8 -3 16 105
use FILL  FILL_1938
timestamp 1714281807
transform 1 0 464 0 1 1570
box -8 -3 16 105
use FILL  FILL_1939
timestamp 1714281807
transform 1 0 456 0 1 1570
box -8 -3 16 105
use FILL  FILL_1940
timestamp 1714281807
transform 1 0 408 0 1 1570
box -8 -3 16 105
use FILL  FILL_1941
timestamp 1714281807
transform 1 0 400 0 1 1570
box -8 -3 16 105
use FILL  FILL_1942
timestamp 1714281807
transform 1 0 392 0 1 1570
box -8 -3 16 105
use FILL  FILL_1943
timestamp 1714281807
transform 1 0 384 0 1 1570
box -8 -3 16 105
use FILL  FILL_1944
timestamp 1714281807
transform 1 0 376 0 1 1570
box -8 -3 16 105
use FILL  FILL_1945
timestamp 1714281807
transform 1 0 368 0 1 1570
box -8 -3 16 105
use FILL  FILL_1946
timestamp 1714281807
transform 1 0 328 0 1 1570
box -8 -3 16 105
use FILL  FILL_1947
timestamp 1714281807
transform 1 0 320 0 1 1570
box -8 -3 16 105
use FILL  FILL_1948
timestamp 1714281807
transform 1 0 312 0 1 1570
box -8 -3 16 105
use FILL  FILL_1949
timestamp 1714281807
transform 1 0 304 0 1 1570
box -8 -3 16 105
use FILL  FILL_1950
timestamp 1714281807
transform 1 0 296 0 1 1570
box -8 -3 16 105
use FILL  FILL_1951
timestamp 1714281807
transform 1 0 288 0 1 1570
box -8 -3 16 105
use FILL  FILL_1952
timestamp 1714281807
transform 1 0 280 0 1 1570
box -8 -3 16 105
use FILL  FILL_1953
timestamp 1714281807
transform 1 0 248 0 1 1570
box -8 -3 16 105
use FILL  FILL_1954
timestamp 1714281807
transform 1 0 240 0 1 1570
box -8 -3 16 105
use FILL  FILL_1955
timestamp 1714281807
transform 1 0 232 0 1 1570
box -8 -3 16 105
use FILL  FILL_1956
timestamp 1714281807
transform 1 0 224 0 1 1570
box -8 -3 16 105
use FILL  FILL_1957
timestamp 1714281807
transform 1 0 216 0 1 1570
box -8 -3 16 105
use FILL  FILL_1958
timestamp 1714281807
transform 1 0 208 0 1 1570
box -8 -3 16 105
use FILL  FILL_1959
timestamp 1714281807
transform 1 0 184 0 1 1570
box -8 -3 16 105
use FILL  FILL_1960
timestamp 1714281807
transform 1 0 176 0 1 1570
box -8 -3 16 105
use FILL  FILL_1961
timestamp 1714281807
transform 1 0 168 0 1 1570
box -8 -3 16 105
use FILL  FILL_1962
timestamp 1714281807
transform 1 0 160 0 1 1570
box -8 -3 16 105
use FILL  FILL_1963
timestamp 1714281807
transform 1 0 152 0 1 1570
box -8 -3 16 105
use FILL  FILL_1964
timestamp 1714281807
transform 1 0 144 0 1 1570
box -8 -3 16 105
use FILL  FILL_1965
timestamp 1714281807
transform 1 0 136 0 1 1570
box -8 -3 16 105
use FILL  FILL_1966
timestamp 1714281807
transform 1 0 128 0 1 1570
box -8 -3 16 105
use FILL  FILL_1967
timestamp 1714281807
transform 1 0 120 0 1 1570
box -8 -3 16 105
use FILL  FILL_1968
timestamp 1714281807
transform 1 0 112 0 1 1570
box -8 -3 16 105
use FILL  FILL_1969
timestamp 1714281807
transform 1 0 104 0 1 1570
box -8 -3 16 105
use FILL  FILL_1970
timestamp 1714281807
transform 1 0 96 0 1 1570
box -8 -3 16 105
use FILL  FILL_1971
timestamp 1714281807
transform 1 0 88 0 1 1570
box -8 -3 16 105
use FILL  FILL_1972
timestamp 1714281807
transform 1 0 80 0 1 1570
box -8 -3 16 105
use FILL  FILL_1973
timestamp 1714281807
transform 1 0 72 0 1 1570
box -8 -3 16 105
use FILL  FILL_1974
timestamp 1714281807
transform 1 0 3000 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1975
timestamp 1714281807
transform 1 0 2992 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1976
timestamp 1714281807
transform 1 0 2984 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1977
timestamp 1714281807
transform 1 0 2976 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1978
timestamp 1714281807
transform 1 0 2968 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1979
timestamp 1714281807
transform 1 0 2960 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1980
timestamp 1714281807
transform 1 0 2952 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1981
timestamp 1714281807
transform 1 0 2944 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1982
timestamp 1714281807
transform 1 0 2936 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1983
timestamp 1714281807
transform 1 0 2928 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1984
timestamp 1714281807
transform 1 0 2920 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1985
timestamp 1714281807
transform 1 0 2912 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1986
timestamp 1714281807
transform 1 0 2904 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1987
timestamp 1714281807
transform 1 0 2896 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1988
timestamp 1714281807
transform 1 0 2888 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1989
timestamp 1714281807
transform 1 0 2880 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1990
timestamp 1714281807
transform 1 0 2872 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1991
timestamp 1714281807
transform 1 0 2768 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1992
timestamp 1714281807
transform 1 0 2760 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1993
timestamp 1714281807
transform 1 0 2752 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1994
timestamp 1714281807
transform 1 0 2744 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1995
timestamp 1714281807
transform 1 0 2736 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1996
timestamp 1714281807
transform 1 0 2704 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1997
timestamp 1714281807
transform 1 0 2696 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1998
timestamp 1714281807
transform 1 0 2688 0 -1 1570
box -8 -3 16 105
use FILL  FILL_1999
timestamp 1714281807
transform 1 0 2664 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2000
timestamp 1714281807
transform 1 0 2656 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2001
timestamp 1714281807
transform 1 0 2648 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2002
timestamp 1714281807
transform 1 0 2640 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2003
timestamp 1714281807
transform 1 0 2600 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2004
timestamp 1714281807
transform 1 0 2592 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2005
timestamp 1714281807
transform 1 0 2584 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2006
timestamp 1714281807
transform 1 0 2576 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2007
timestamp 1714281807
transform 1 0 2568 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2008
timestamp 1714281807
transform 1 0 2560 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2009
timestamp 1714281807
transform 1 0 2536 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2010
timestamp 1714281807
transform 1 0 2528 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2011
timestamp 1714281807
transform 1 0 2520 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2012
timestamp 1714281807
transform 1 0 2480 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2013
timestamp 1714281807
transform 1 0 2472 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2014
timestamp 1714281807
transform 1 0 2464 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2015
timestamp 1714281807
transform 1 0 2456 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2016
timestamp 1714281807
transform 1 0 2448 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2017
timestamp 1714281807
transform 1 0 2440 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2018
timestamp 1714281807
transform 1 0 2432 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2019
timestamp 1714281807
transform 1 0 2400 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2020
timestamp 1714281807
transform 1 0 2392 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2021
timestamp 1714281807
transform 1 0 2384 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2022
timestamp 1714281807
transform 1 0 2376 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2023
timestamp 1714281807
transform 1 0 2272 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2024
timestamp 1714281807
transform 1 0 2264 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2025
timestamp 1714281807
transform 1 0 2160 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2026
timestamp 1714281807
transform 1 0 2152 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2027
timestamp 1714281807
transform 1 0 2144 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2028
timestamp 1714281807
transform 1 0 2136 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2029
timestamp 1714281807
transform 1 0 2072 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2030
timestamp 1714281807
transform 1 0 2064 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2031
timestamp 1714281807
transform 1 0 2056 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2032
timestamp 1714281807
transform 1 0 1952 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2033
timestamp 1714281807
transform 1 0 1848 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2034
timestamp 1714281807
transform 1 0 1840 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2035
timestamp 1714281807
transform 1 0 1712 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2036
timestamp 1714281807
transform 1 0 1704 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2037
timestamp 1714281807
transform 1 0 1696 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2038
timestamp 1714281807
transform 1 0 1688 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2039
timestamp 1714281807
transform 1 0 1640 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2040
timestamp 1714281807
transform 1 0 1632 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2041
timestamp 1714281807
transform 1 0 1624 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2042
timestamp 1714281807
transform 1 0 1616 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2043
timestamp 1714281807
transform 1 0 1608 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2044
timestamp 1714281807
transform 1 0 1600 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2045
timestamp 1714281807
transform 1 0 1592 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2046
timestamp 1714281807
transform 1 0 1552 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2047
timestamp 1714281807
transform 1 0 1528 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2048
timestamp 1714281807
transform 1 0 1520 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2049
timestamp 1714281807
transform 1 0 1512 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2050
timestamp 1714281807
transform 1 0 1504 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2051
timestamp 1714281807
transform 1 0 1496 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2052
timestamp 1714281807
transform 1 0 1488 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2053
timestamp 1714281807
transform 1 0 1480 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2054
timestamp 1714281807
transform 1 0 1448 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2055
timestamp 1714281807
transform 1 0 1440 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2056
timestamp 1714281807
transform 1 0 1432 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2057
timestamp 1714281807
transform 1 0 1424 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2058
timestamp 1714281807
transform 1 0 1416 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2059
timestamp 1714281807
transform 1 0 1408 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2060
timestamp 1714281807
transform 1 0 1400 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2061
timestamp 1714281807
transform 1 0 1392 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2062
timestamp 1714281807
transform 1 0 1344 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2063
timestamp 1714281807
transform 1 0 1336 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2064
timestamp 1714281807
transform 1 0 1328 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2065
timestamp 1714281807
transform 1 0 1320 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2066
timestamp 1714281807
transform 1 0 1312 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2067
timestamp 1714281807
transform 1 0 1288 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2068
timestamp 1714281807
transform 1 0 1280 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2069
timestamp 1714281807
transform 1 0 1272 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2070
timestamp 1714281807
transform 1 0 1264 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2071
timestamp 1714281807
transform 1 0 1256 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2072
timestamp 1714281807
transform 1 0 1208 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2073
timestamp 1714281807
transform 1 0 1200 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2074
timestamp 1714281807
transform 1 0 1192 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2075
timestamp 1714281807
transform 1 0 1184 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2076
timestamp 1714281807
transform 1 0 1176 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2077
timestamp 1714281807
transform 1 0 1168 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2078
timestamp 1714281807
transform 1 0 1160 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2079
timestamp 1714281807
transform 1 0 1112 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2080
timestamp 1714281807
transform 1 0 1104 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2081
timestamp 1714281807
transform 1 0 1096 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2082
timestamp 1714281807
transform 1 0 1088 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2083
timestamp 1714281807
transform 1 0 1080 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2084
timestamp 1714281807
transform 1 0 1072 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2085
timestamp 1714281807
transform 1 0 1064 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2086
timestamp 1714281807
transform 1 0 1056 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2087
timestamp 1714281807
transform 1 0 1008 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2088
timestamp 1714281807
transform 1 0 1000 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2089
timestamp 1714281807
transform 1 0 992 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2090
timestamp 1714281807
transform 1 0 984 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2091
timestamp 1714281807
transform 1 0 976 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2092
timestamp 1714281807
transform 1 0 968 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2093
timestamp 1714281807
transform 1 0 960 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2094
timestamp 1714281807
transform 1 0 952 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2095
timestamp 1714281807
transform 1 0 896 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2096
timestamp 1714281807
transform 1 0 888 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2097
timestamp 1714281807
transform 1 0 880 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2098
timestamp 1714281807
transform 1 0 776 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2099
timestamp 1714281807
transform 1 0 768 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2100
timestamp 1714281807
transform 1 0 760 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2101
timestamp 1714281807
transform 1 0 752 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2102
timestamp 1714281807
transform 1 0 744 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2103
timestamp 1714281807
transform 1 0 712 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2104
timestamp 1714281807
transform 1 0 704 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2105
timestamp 1714281807
transform 1 0 696 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2106
timestamp 1714281807
transform 1 0 688 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2107
timestamp 1714281807
transform 1 0 656 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2108
timestamp 1714281807
transform 1 0 648 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2109
timestamp 1714281807
transform 1 0 640 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2110
timestamp 1714281807
transform 1 0 632 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2111
timestamp 1714281807
transform 1 0 624 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2112
timestamp 1714281807
transform 1 0 616 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2113
timestamp 1714281807
transform 1 0 608 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2114
timestamp 1714281807
transform 1 0 568 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2115
timestamp 1714281807
transform 1 0 560 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2116
timestamp 1714281807
transform 1 0 552 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2117
timestamp 1714281807
transform 1 0 544 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2118
timestamp 1714281807
transform 1 0 520 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2119
timestamp 1714281807
transform 1 0 512 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2120
timestamp 1714281807
transform 1 0 504 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2121
timestamp 1714281807
transform 1 0 496 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2122
timestamp 1714281807
transform 1 0 488 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2123
timestamp 1714281807
transform 1 0 456 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2124
timestamp 1714281807
transform 1 0 448 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2125
timestamp 1714281807
transform 1 0 440 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2126
timestamp 1714281807
transform 1 0 432 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2127
timestamp 1714281807
transform 1 0 424 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2128
timestamp 1714281807
transform 1 0 416 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2129
timestamp 1714281807
transform 1 0 384 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2130
timestamp 1714281807
transform 1 0 376 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2131
timestamp 1714281807
transform 1 0 368 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2132
timestamp 1714281807
transform 1 0 360 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2133
timestamp 1714281807
transform 1 0 352 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2134
timestamp 1714281807
transform 1 0 328 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2135
timestamp 1714281807
transform 1 0 320 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2136
timestamp 1714281807
transform 1 0 312 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2137
timestamp 1714281807
transform 1 0 304 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2138
timestamp 1714281807
transform 1 0 296 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2139
timestamp 1714281807
transform 1 0 248 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2140
timestamp 1714281807
transform 1 0 240 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2141
timestamp 1714281807
transform 1 0 232 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2142
timestamp 1714281807
transform 1 0 224 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2143
timestamp 1714281807
transform 1 0 216 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2144
timestamp 1714281807
transform 1 0 112 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2145
timestamp 1714281807
transform 1 0 104 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2146
timestamp 1714281807
transform 1 0 96 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2147
timestamp 1714281807
transform 1 0 88 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2148
timestamp 1714281807
transform 1 0 80 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2149
timestamp 1714281807
transform 1 0 72 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2150
timestamp 1714281807
transform 1 0 3000 0 1 1370
box -8 -3 16 105
use FILL  FILL_2151
timestamp 1714281807
transform 1 0 2992 0 1 1370
box -8 -3 16 105
use FILL  FILL_2152
timestamp 1714281807
transform 1 0 2984 0 1 1370
box -8 -3 16 105
use FILL  FILL_2153
timestamp 1714281807
transform 1 0 2880 0 1 1370
box -8 -3 16 105
use FILL  FILL_2154
timestamp 1714281807
transform 1 0 2872 0 1 1370
box -8 -3 16 105
use FILL  FILL_2155
timestamp 1714281807
transform 1 0 2864 0 1 1370
box -8 -3 16 105
use FILL  FILL_2156
timestamp 1714281807
transform 1 0 2824 0 1 1370
box -8 -3 16 105
use FILL  FILL_2157
timestamp 1714281807
transform 1 0 2816 0 1 1370
box -8 -3 16 105
use FILL  FILL_2158
timestamp 1714281807
transform 1 0 2808 0 1 1370
box -8 -3 16 105
use FILL  FILL_2159
timestamp 1714281807
transform 1 0 2800 0 1 1370
box -8 -3 16 105
use FILL  FILL_2160
timestamp 1714281807
transform 1 0 2792 0 1 1370
box -8 -3 16 105
use FILL  FILL_2161
timestamp 1714281807
transform 1 0 2784 0 1 1370
box -8 -3 16 105
use FILL  FILL_2162
timestamp 1714281807
transform 1 0 2776 0 1 1370
box -8 -3 16 105
use FILL  FILL_2163
timestamp 1714281807
transform 1 0 2728 0 1 1370
box -8 -3 16 105
use FILL  FILL_2164
timestamp 1714281807
transform 1 0 2720 0 1 1370
box -8 -3 16 105
use FILL  FILL_2165
timestamp 1714281807
transform 1 0 2712 0 1 1370
box -8 -3 16 105
use FILL  FILL_2166
timestamp 1714281807
transform 1 0 2704 0 1 1370
box -8 -3 16 105
use FILL  FILL_2167
timestamp 1714281807
transform 1 0 2696 0 1 1370
box -8 -3 16 105
use FILL  FILL_2168
timestamp 1714281807
transform 1 0 2592 0 1 1370
box -8 -3 16 105
use FILL  FILL_2169
timestamp 1714281807
transform 1 0 2584 0 1 1370
box -8 -3 16 105
use FILL  FILL_2170
timestamp 1714281807
transform 1 0 2480 0 1 1370
box -8 -3 16 105
use FILL  FILL_2171
timestamp 1714281807
transform 1 0 2376 0 1 1370
box -8 -3 16 105
use FILL  FILL_2172
timestamp 1714281807
transform 1 0 2368 0 1 1370
box -8 -3 16 105
use FILL  FILL_2173
timestamp 1714281807
transform 1 0 2360 0 1 1370
box -8 -3 16 105
use FILL  FILL_2174
timestamp 1714281807
transform 1 0 2336 0 1 1370
box -8 -3 16 105
use FILL  FILL_2175
timestamp 1714281807
transform 1 0 2328 0 1 1370
box -8 -3 16 105
use FILL  FILL_2176
timestamp 1714281807
transform 1 0 2320 0 1 1370
box -8 -3 16 105
use FILL  FILL_2177
timestamp 1714281807
transform 1 0 2312 0 1 1370
box -8 -3 16 105
use FILL  FILL_2178
timestamp 1714281807
transform 1 0 2304 0 1 1370
box -8 -3 16 105
use FILL  FILL_2179
timestamp 1714281807
transform 1 0 2296 0 1 1370
box -8 -3 16 105
use FILL  FILL_2180
timestamp 1714281807
transform 1 0 2288 0 1 1370
box -8 -3 16 105
use FILL  FILL_2181
timestamp 1714281807
transform 1 0 2280 0 1 1370
box -8 -3 16 105
use FILL  FILL_2182
timestamp 1714281807
transform 1 0 2272 0 1 1370
box -8 -3 16 105
use FILL  FILL_2183
timestamp 1714281807
transform 1 0 2264 0 1 1370
box -8 -3 16 105
use FILL  FILL_2184
timestamp 1714281807
transform 1 0 2160 0 1 1370
box -8 -3 16 105
use FILL  FILL_2185
timestamp 1714281807
transform 1 0 2152 0 1 1370
box -8 -3 16 105
use FILL  FILL_2186
timestamp 1714281807
transform 1 0 2144 0 1 1370
box -8 -3 16 105
use FILL  FILL_2187
timestamp 1714281807
transform 1 0 2136 0 1 1370
box -8 -3 16 105
use FILL  FILL_2188
timestamp 1714281807
transform 1 0 2104 0 1 1370
box -8 -3 16 105
use FILL  FILL_2189
timestamp 1714281807
transform 1 0 2096 0 1 1370
box -8 -3 16 105
use FILL  FILL_2190
timestamp 1714281807
transform 1 0 2088 0 1 1370
box -8 -3 16 105
use FILL  FILL_2191
timestamp 1714281807
transform 1 0 2064 0 1 1370
box -8 -3 16 105
use FILL  FILL_2192
timestamp 1714281807
transform 1 0 2056 0 1 1370
box -8 -3 16 105
use FILL  FILL_2193
timestamp 1714281807
transform 1 0 2048 0 1 1370
box -8 -3 16 105
use FILL  FILL_2194
timestamp 1714281807
transform 1 0 2040 0 1 1370
box -8 -3 16 105
use FILL  FILL_2195
timestamp 1714281807
transform 1 0 1976 0 1 1370
box -8 -3 16 105
use FILL  FILL_2196
timestamp 1714281807
transform 1 0 1968 0 1 1370
box -8 -3 16 105
use FILL  FILL_2197
timestamp 1714281807
transform 1 0 1960 0 1 1370
box -8 -3 16 105
use FILL  FILL_2198
timestamp 1714281807
transform 1 0 1856 0 1 1370
box -8 -3 16 105
use FILL  FILL_2199
timestamp 1714281807
transform 1 0 1848 0 1 1370
box -8 -3 16 105
use FILL  FILL_2200
timestamp 1714281807
transform 1 0 1840 0 1 1370
box -8 -3 16 105
use FILL  FILL_2201
timestamp 1714281807
transform 1 0 1832 0 1 1370
box -8 -3 16 105
use FILL  FILL_2202
timestamp 1714281807
transform 1 0 1784 0 1 1370
box -8 -3 16 105
use FILL  FILL_2203
timestamp 1714281807
transform 1 0 1776 0 1 1370
box -8 -3 16 105
use FILL  FILL_2204
timestamp 1714281807
transform 1 0 1768 0 1 1370
box -8 -3 16 105
use FILL  FILL_2205
timestamp 1714281807
transform 1 0 1760 0 1 1370
box -8 -3 16 105
use FILL  FILL_2206
timestamp 1714281807
transform 1 0 1752 0 1 1370
box -8 -3 16 105
use FILL  FILL_2207
timestamp 1714281807
transform 1 0 1568 0 1 1370
box -8 -3 16 105
use FILL  FILL_2208
timestamp 1714281807
transform 1 0 1560 0 1 1370
box -8 -3 16 105
use FILL  FILL_2209
timestamp 1714281807
transform 1 0 1528 0 1 1370
box -8 -3 16 105
use FILL  FILL_2210
timestamp 1714281807
transform 1 0 1520 0 1 1370
box -8 -3 16 105
use FILL  FILL_2211
timestamp 1714281807
transform 1 0 1512 0 1 1370
box -8 -3 16 105
use FILL  FILL_2212
timestamp 1714281807
transform 1 0 1504 0 1 1370
box -8 -3 16 105
use FILL  FILL_2213
timestamp 1714281807
transform 1 0 1472 0 1 1370
box -8 -3 16 105
use FILL  FILL_2214
timestamp 1714281807
transform 1 0 1464 0 1 1370
box -8 -3 16 105
use FILL  FILL_2215
timestamp 1714281807
transform 1 0 1456 0 1 1370
box -8 -3 16 105
use FILL  FILL_2216
timestamp 1714281807
transform 1 0 1448 0 1 1370
box -8 -3 16 105
use FILL  FILL_2217
timestamp 1714281807
transform 1 0 1440 0 1 1370
box -8 -3 16 105
use FILL  FILL_2218
timestamp 1714281807
transform 1 0 1408 0 1 1370
box -8 -3 16 105
use FILL  FILL_2219
timestamp 1714281807
transform 1 0 1400 0 1 1370
box -8 -3 16 105
use FILL  FILL_2220
timestamp 1714281807
transform 1 0 1392 0 1 1370
box -8 -3 16 105
use FILL  FILL_2221
timestamp 1714281807
transform 1 0 1384 0 1 1370
box -8 -3 16 105
use FILL  FILL_2222
timestamp 1714281807
transform 1 0 1352 0 1 1370
box -8 -3 16 105
use FILL  FILL_2223
timestamp 1714281807
transform 1 0 1344 0 1 1370
box -8 -3 16 105
use FILL  FILL_2224
timestamp 1714281807
transform 1 0 1336 0 1 1370
box -8 -3 16 105
use FILL  FILL_2225
timestamp 1714281807
transform 1 0 1328 0 1 1370
box -8 -3 16 105
use FILL  FILL_2226
timestamp 1714281807
transform 1 0 1320 0 1 1370
box -8 -3 16 105
use FILL  FILL_2227
timestamp 1714281807
transform 1 0 1312 0 1 1370
box -8 -3 16 105
use FILL  FILL_2228
timestamp 1714281807
transform 1 0 1264 0 1 1370
box -8 -3 16 105
use FILL  FILL_2229
timestamp 1714281807
transform 1 0 1256 0 1 1370
box -8 -3 16 105
use FILL  FILL_2230
timestamp 1714281807
transform 1 0 1248 0 1 1370
box -8 -3 16 105
use FILL  FILL_2231
timestamp 1714281807
transform 1 0 1240 0 1 1370
box -8 -3 16 105
use FILL  FILL_2232
timestamp 1714281807
transform 1 0 1232 0 1 1370
box -8 -3 16 105
use FILL  FILL_2233
timestamp 1714281807
transform 1 0 1224 0 1 1370
box -8 -3 16 105
use FILL  FILL_2234
timestamp 1714281807
transform 1 0 1216 0 1 1370
box -8 -3 16 105
use FILL  FILL_2235
timestamp 1714281807
transform 1 0 1176 0 1 1370
box -8 -3 16 105
use FILL  FILL_2236
timestamp 1714281807
transform 1 0 1168 0 1 1370
box -8 -3 16 105
use FILL  FILL_2237
timestamp 1714281807
transform 1 0 1160 0 1 1370
box -8 -3 16 105
use FILL  FILL_2238
timestamp 1714281807
transform 1 0 1152 0 1 1370
box -8 -3 16 105
use FILL  FILL_2239
timestamp 1714281807
transform 1 0 1144 0 1 1370
box -8 -3 16 105
use FILL  FILL_2240
timestamp 1714281807
transform 1 0 1136 0 1 1370
box -8 -3 16 105
use FILL  FILL_2241
timestamp 1714281807
transform 1 0 1128 0 1 1370
box -8 -3 16 105
use FILL  FILL_2242
timestamp 1714281807
transform 1 0 1080 0 1 1370
box -8 -3 16 105
use FILL  FILL_2243
timestamp 1714281807
transform 1 0 1072 0 1 1370
box -8 -3 16 105
use FILL  FILL_2244
timestamp 1714281807
transform 1 0 1064 0 1 1370
box -8 -3 16 105
use FILL  FILL_2245
timestamp 1714281807
transform 1 0 1056 0 1 1370
box -8 -3 16 105
use FILL  FILL_2246
timestamp 1714281807
transform 1 0 1048 0 1 1370
box -8 -3 16 105
use FILL  FILL_2247
timestamp 1714281807
transform 1 0 1024 0 1 1370
box -8 -3 16 105
use FILL  FILL_2248
timestamp 1714281807
transform 1 0 984 0 1 1370
box -8 -3 16 105
use FILL  FILL_2249
timestamp 1714281807
transform 1 0 976 0 1 1370
box -8 -3 16 105
use FILL  FILL_2250
timestamp 1714281807
transform 1 0 968 0 1 1370
box -8 -3 16 105
use FILL  FILL_2251
timestamp 1714281807
transform 1 0 928 0 1 1370
box -8 -3 16 105
use FILL  FILL_2252
timestamp 1714281807
transform 1 0 920 0 1 1370
box -8 -3 16 105
use FILL  FILL_2253
timestamp 1714281807
transform 1 0 912 0 1 1370
box -8 -3 16 105
use FILL  FILL_2254
timestamp 1714281807
transform 1 0 888 0 1 1370
box -8 -3 16 105
use FILL  FILL_2255
timestamp 1714281807
transform 1 0 880 0 1 1370
box -8 -3 16 105
use FILL  FILL_2256
timestamp 1714281807
transform 1 0 872 0 1 1370
box -8 -3 16 105
use FILL  FILL_2257
timestamp 1714281807
transform 1 0 848 0 1 1370
box -8 -3 16 105
use FILL  FILL_2258
timestamp 1714281807
transform 1 0 840 0 1 1370
box -8 -3 16 105
use FILL  FILL_2259
timestamp 1714281807
transform 1 0 808 0 1 1370
box -8 -3 16 105
use FILL  FILL_2260
timestamp 1714281807
transform 1 0 800 0 1 1370
box -8 -3 16 105
use FILL  FILL_2261
timestamp 1714281807
transform 1 0 792 0 1 1370
box -8 -3 16 105
use FILL  FILL_2262
timestamp 1714281807
transform 1 0 784 0 1 1370
box -8 -3 16 105
use FILL  FILL_2263
timestamp 1714281807
transform 1 0 776 0 1 1370
box -8 -3 16 105
use FILL  FILL_2264
timestamp 1714281807
transform 1 0 736 0 1 1370
box -8 -3 16 105
use FILL  FILL_2265
timestamp 1714281807
transform 1 0 728 0 1 1370
box -8 -3 16 105
use FILL  FILL_2266
timestamp 1714281807
transform 1 0 720 0 1 1370
box -8 -3 16 105
use FILL  FILL_2267
timestamp 1714281807
transform 1 0 712 0 1 1370
box -8 -3 16 105
use FILL  FILL_2268
timestamp 1714281807
transform 1 0 704 0 1 1370
box -8 -3 16 105
use FILL  FILL_2269
timestamp 1714281807
transform 1 0 656 0 1 1370
box -8 -3 16 105
use FILL  FILL_2270
timestamp 1714281807
transform 1 0 648 0 1 1370
box -8 -3 16 105
use FILL  FILL_2271
timestamp 1714281807
transform 1 0 640 0 1 1370
box -8 -3 16 105
use FILL  FILL_2272
timestamp 1714281807
transform 1 0 536 0 1 1370
box -8 -3 16 105
use FILL  FILL_2273
timestamp 1714281807
transform 1 0 528 0 1 1370
box -8 -3 16 105
use FILL  FILL_2274
timestamp 1714281807
transform 1 0 520 0 1 1370
box -8 -3 16 105
use FILL  FILL_2275
timestamp 1714281807
transform 1 0 512 0 1 1370
box -8 -3 16 105
use FILL  FILL_2276
timestamp 1714281807
transform 1 0 504 0 1 1370
box -8 -3 16 105
use FILL  FILL_2277
timestamp 1714281807
transform 1 0 472 0 1 1370
box -8 -3 16 105
use FILL  FILL_2278
timestamp 1714281807
transform 1 0 464 0 1 1370
box -8 -3 16 105
use FILL  FILL_2279
timestamp 1714281807
transform 1 0 440 0 1 1370
box -8 -3 16 105
use FILL  FILL_2280
timestamp 1714281807
transform 1 0 432 0 1 1370
box -8 -3 16 105
use FILL  FILL_2281
timestamp 1714281807
transform 1 0 424 0 1 1370
box -8 -3 16 105
use FILL  FILL_2282
timestamp 1714281807
transform 1 0 416 0 1 1370
box -8 -3 16 105
use FILL  FILL_2283
timestamp 1714281807
transform 1 0 384 0 1 1370
box -8 -3 16 105
use FILL  FILL_2284
timestamp 1714281807
transform 1 0 376 0 1 1370
box -8 -3 16 105
use FILL  FILL_2285
timestamp 1714281807
transform 1 0 368 0 1 1370
box -8 -3 16 105
use FILL  FILL_2286
timestamp 1714281807
transform 1 0 360 0 1 1370
box -8 -3 16 105
use FILL  FILL_2287
timestamp 1714281807
transform 1 0 352 0 1 1370
box -8 -3 16 105
use FILL  FILL_2288
timestamp 1714281807
transform 1 0 344 0 1 1370
box -8 -3 16 105
use FILL  FILL_2289
timestamp 1714281807
transform 1 0 304 0 1 1370
box -8 -3 16 105
use FILL  FILL_2290
timestamp 1714281807
transform 1 0 296 0 1 1370
box -8 -3 16 105
use FILL  FILL_2291
timestamp 1714281807
transform 1 0 288 0 1 1370
box -8 -3 16 105
use FILL  FILL_2292
timestamp 1714281807
transform 1 0 280 0 1 1370
box -8 -3 16 105
use FILL  FILL_2293
timestamp 1714281807
transform 1 0 272 0 1 1370
box -8 -3 16 105
use FILL  FILL_2294
timestamp 1714281807
transform 1 0 240 0 1 1370
box -8 -3 16 105
use FILL  FILL_2295
timestamp 1714281807
transform 1 0 232 0 1 1370
box -8 -3 16 105
use FILL  FILL_2296
timestamp 1714281807
transform 1 0 224 0 1 1370
box -8 -3 16 105
use FILL  FILL_2297
timestamp 1714281807
transform 1 0 120 0 1 1370
box -8 -3 16 105
use FILL  FILL_2298
timestamp 1714281807
transform 1 0 112 0 1 1370
box -8 -3 16 105
use FILL  FILL_2299
timestamp 1714281807
transform 1 0 104 0 1 1370
box -8 -3 16 105
use FILL  FILL_2300
timestamp 1714281807
transform 1 0 96 0 1 1370
box -8 -3 16 105
use FILL  FILL_2301
timestamp 1714281807
transform 1 0 88 0 1 1370
box -8 -3 16 105
use FILL  FILL_2302
timestamp 1714281807
transform 1 0 80 0 1 1370
box -8 -3 16 105
use FILL  FILL_2303
timestamp 1714281807
transform 1 0 72 0 1 1370
box -8 -3 16 105
use FILL  FILL_2304
timestamp 1714281807
transform 1 0 3000 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2305
timestamp 1714281807
transform 1 0 2992 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2306
timestamp 1714281807
transform 1 0 2984 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2307
timestamp 1714281807
transform 1 0 2976 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2308
timestamp 1714281807
transform 1 0 2968 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2309
timestamp 1714281807
transform 1 0 2960 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2310
timestamp 1714281807
transform 1 0 2952 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2311
timestamp 1714281807
transform 1 0 2944 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2312
timestamp 1714281807
transform 1 0 2936 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2313
timestamp 1714281807
transform 1 0 2912 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2314
timestamp 1714281807
transform 1 0 2904 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2315
timestamp 1714281807
transform 1 0 2784 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2316
timestamp 1714281807
transform 1 0 2776 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2317
timestamp 1714281807
transform 1 0 2736 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2318
timestamp 1714281807
transform 1 0 2728 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2319
timestamp 1714281807
transform 1 0 2664 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2320
timestamp 1714281807
transform 1 0 2656 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2321
timestamp 1714281807
transform 1 0 2616 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2322
timestamp 1714281807
transform 1 0 2608 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2323
timestamp 1714281807
transform 1 0 2600 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2324
timestamp 1714281807
transform 1 0 2592 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2325
timestamp 1714281807
transform 1 0 2584 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2326
timestamp 1714281807
transform 1 0 2536 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2327
timestamp 1714281807
transform 1 0 2528 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2328
timestamp 1714281807
transform 1 0 2520 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2329
timestamp 1714281807
transform 1 0 2512 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2330
timestamp 1714281807
transform 1 0 2504 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2331
timestamp 1714281807
transform 1 0 2496 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2332
timestamp 1714281807
transform 1 0 2464 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2333
timestamp 1714281807
transform 1 0 2456 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2334
timestamp 1714281807
transform 1 0 2448 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2335
timestamp 1714281807
transform 1 0 2408 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2336
timestamp 1714281807
transform 1 0 2400 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2337
timestamp 1714281807
transform 1 0 2392 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2338
timestamp 1714281807
transform 1 0 2384 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2339
timestamp 1714281807
transform 1 0 2376 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2340
timestamp 1714281807
transform 1 0 2368 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2341
timestamp 1714281807
transform 1 0 2360 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2342
timestamp 1714281807
transform 1 0 2304 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2343
timestamp 1714281807
transform 1 0 2296 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2344
timestamp 1714281807
transform 1 0 2192 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2345
timestamp 1714281807
transform 1 0 2184 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2346
timestamp 1714281807
transform 1 0 2176 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2347
timestamp 1714281807
transform 1 0 2096 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2348
timestamp 1714281807
transform 1 0 2088 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2349
timestamp 1714281807
transform 1 0 2080 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2350
timestamp 1714281807
transform 1 0 2072 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2351
timestamp 1714281807
transform 1 0 2064 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2352
timestamp 1714281807
transform 1 0 2056 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2353
timestamp 1714281807
transform 1 0 2048 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2354
timestamp 1714281807
transform 1 0 1992 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2355
timestamp 1714281807
transform 1 0 1984 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2356
timestamp 1714281807
transform 1 0 1880 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2357
timestamp 1714281807
transform 1 0 1872 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2358
timestamp 1714281807
transform 1 0 1864 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2359
timestamp 1714281807
transform 1 0 1824 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2360
timestamp 1714281807
transform 1 0 1816 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2361
timestamp 1714281807
transform 1 0 1808 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2362
timestamp 1714281807
transform 1 0 1800 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2363
timestamp 1714281807
transform 1 0 1752 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2364
timestamp 1714281807
transform 1 0 1744 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2365
timestamp 1714281807
transform 1 0 1736 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2366
timestamp 1714281807
transform 1 0 1728 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2367
timestamp 1714281807
transform 1 0 1664 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2368
timestamp 1714281807
transform 1 0 1632 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2369
timestamp 1714281807
transform 1 0 1624 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2370
timestamp 1714281807
transform 1 0 1616 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2371
timestamp 1714281807
transform 1 0 1608 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2372
timestamp 1714281807
transform 1 0 1600 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2373
timestamp 1714281807
transform 1 0 1592 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2374
timestamp 1714281807
transform 1 0 1584 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2375
timestamp 1714281807
transform 1 0 1544 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2376
timestamp 1714281807
transform 1 0 1536 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2377
timestamp 1714281807
transform 1 0 1528 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2378
timestamp 1714281807
transform 1 0 1520 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2379
timestamp 1714281807
transform 1 0 1512 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2380
timestamp 1714281807
transform 1 0 1504 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2381
timestamp 1714281807
transform 1 0 1496 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2382
timestamp 1714281807
transform 1 0 1464 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2383
timestamp 1714281807
transform 1 0 1456 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2384
timestamp 1714281807
transform 1 0 1448 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2385
timestamp 1714281807
transform 1 0 1440 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2386
timestamp 1714281807
transform 1 0 1432 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2387
timestamp 1714281807
transform 1 0 1408 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2388
timestamp 1714281807
transform 1 0 1400 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2389
timestamp 1714281807
transform 1 0 1368 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2390
timestamp 1714281807
transform 1 0 1312 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2391
timestamp 1714281807
transform 1 0 1304 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2392
timestamp 1714281807
transform 1 0 1296 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2393
timestamp 1714281807
transform 1 0 1264 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2394
timestamp 1714281807
transform 1 0 1216 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2395
timestamp 1714281807
transform 1 0 1208 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2396
timestamp 1714281807
transform 1 0 1200 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2397
timestamp 1714281807
transform 1 0 1192 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2398
timestamp 1714281807
transform 1 0 1184 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2399
timestamp 1714281807
transform 1 0 1136 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2400
timestamp 1714281807
transform 1 0 1128 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2401
timestamp 1714281807
transform 1 0 1120 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2402
timestamp 1714281807
transform 1 0 1112 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2403
timestamp 1714281807
transform 1 0 1104 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2404
timestamp 1714281807
transform 1 0 1096 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2405
timestamp 1714281807
transform 1 0 1088 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2406
timestamp 1714281807
transform 1 0 1056 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2407
timestamp 1714281807
transform 1 0 1048 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2408
timestamp 1714281807
transform 1 0 1040 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2409
timestamp 1714281807
transform 1 0 1032 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2410
timestamp 1714281807
transform 1 0 1024 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2411
timestamp 1714281807
transform 1 0 1016 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2412
timestamp 1714281807
transform 1 0 960 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2413
timestamp 1714281807
transform 1 0 952 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2414
timestamp 1714281807
transform 1 0 944 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2415
timestamp 1714281807
transform 1 0 936 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2416
timestamp 1714281807
transform 1 0 928 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2417
timestamp 1714281807
transform 1 0 856 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2418
timestamp 1714281807
transform 1 0 848 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2419
timestamp 1714281807
transform 1 0 840 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2420
timestamp 1714281807
transform 1 0 832 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2421
timestamp 1714281807
transform 1 0 824 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2422
timestamp 1714281807
transform 1 0 816 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2423
timestamp 1714281807
transform 1 0 768 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2424
timestamp 1714281807
transform 1 0 760 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2425
timestamp 1714281807
transform 1 0 752 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2426
timestamp 1714281807
transform 1 0 744 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2427
timestamp 1714281807
transform 1 0 736 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2428
timestamp 1714281807
transform 1 0 712 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2429
timestamp 1714281807
transform 1 0 704 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2430
timestamp 1714281807
transform 1 0 696 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2431
timestamp 1714281807
transform 1 0 688 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2432
timestamp 1714281807
transform 1 0 656 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2433
timestamp 1714281807
transform 1 0 648 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2434
timestamp 1714281807
transform 1 0 640 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2435
timestamp 1714281807
transform 1 0 632 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2436
timestamp 1714281807
transform 1 0 528 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2437
timestamp 1714281807
transform 1 0 520 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2438
timestamp 1714281807
transform 1 0 416 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2439
timestamp 1714281807
transform 1 0 408 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2440
timestamp 1714281807
transform 1 0 400 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2441
timestamp 1714281807
transform 1 0 376 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2442
timestamp 1714281807
transform 1 0 368 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2443
timestamp 1714281807
transform 1 0 360 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2444
timestamp 1714281807
transform 1 0 352 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2445
timestamp 1714281807
transform 1 0 328 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2446
timestamp 1714281807
transform 1 0 320 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2447
timestamp 1714281807
transform 1 0 312 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2448
timestamp 1714281807
transform 1 0 208 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2449
timestamp 1714281807
transform 1 0 200 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2450
timestamp 1714281807
transform 1 0 192 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2451
timestamp 1714281807
transform 1 0 184 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2452
timestamp 1714281807
transform 1 0 176 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2453
timestamp 1714281807
transform 1 0 168 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2454
timestamp 1714281807
transform 1 0 160 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2455
timestamp 1714281807
transform 1 0 152 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2456
timestamp 1714281807
transform 1 0 144 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2457
timestamp 1714281807
transform 1 0 136 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2458
timestamp 1714281807
transform 1 0 128 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2459
timestamp 1714281807
transform 1 0 120 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2460
timestamp 1714281807
transform 1 0 112 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2461
timestamp 1714281807
transform 1 0 104 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2462
timestamp 1714281807
transform 1 0 96 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2463
timestamp 1714281807
transform 1 0 88 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2464
timestamp 1714281807
transform 1 0 80 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2465
timestamp 1714281807
transform 1 0 72 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2466
timestamp 1714281807
transform 1 0 3000 0 1 1170
box -8 -3 16 105
use FILL  FILL_2467
timestamp 1714281807
transform 1 0 2896 0 1 1170
box -8 -3 16 105
use FILL  FILL_2468
timestamp 1714281807
transform 1 0 2888 0 1 1170
box -8 -3 16 105
use FILL  FILL_2469
timestamp 1714281807
transform 1 0 2864 0 1 1170
box -8 -3 16 105
use FILL  FILL_2470
timestamp 1714281807
transform 1 0 2856 0 1 1170
box -8 -3 16 105
use FILL  FILL_2471
timestamp 1714281807
transform 1 0 2816 0 1 1170
box -8 -3 16 105
use FILL  FILL_2472
timestamp 1714281807
transform 1 0 2808 0 1 1170
box -8 -3 16 105
use FILL  FILL_2473
timestamp 1714281807
transform 1 0 2800 0 1 1170
box -8 -3 16 105
use FILL  FILL_2474
timestamp 1714281807
transform 1 0 2792 0 1 1170
box -8 -3 16 105
use FILL  FILL_2475
timestamp 1714281807
transform 1 0 2784 0 1 1170
box -8 -3 16 105
use FILL  FILL_2476
timestamp 1714281807
transform 1 0 2776 0 1 1170
box -8 -3 16 105
use FILL  FILL_2477
timestamp 1714281807
transform 1 0 2728 0 1 1170
box -8 -3 16 105
use FILL  FILL_2478
timestamp 1714281807
transform 1 0 2720 0 1 1170
box -8 -3 16 105
use FILL  FILL_2479
timestamp 1714281807
transform 1 0 2712 0 1 1170
box -8 -3 16 105
use FILL  FILL_2480
timestamp 1714281807
transform 1 0 2704 0 1 1170
box -8 -3 16 105
use FILL  FILL_2481
timestamp 1714281807
transform 1 0 2696 0 1 1170
box -8 -3 16 105
use FILL  FILL_2482
timestamp 1714281807
transform 1 0 2576 0 1 1170
box -8 -3 16 105
use FILL  FILL_2483
timestamp 1714281807
transform 1 0 2536 0 1 1170
box -8 -3 16 105
use FILL  FILL_2484
timestamp 1714281807
transform 1 0 2528 0 1 1170
box -8 -3 16 105
use FILL  FILL_2485
timestamp 1714281807
transform 1 0 2496 0 1 1170
box -8 -3 16 105
use FILL  FILL_2486
timestamp 1714281807
transform 1 0 2488 0 1 1170
box -8 -3 16 105
use FILL  FILL_2487
timestamp 1714281807
transform 1 0 2480 0 1 1170
box -8 -3 16 105
use FILL  FILL_2488
timestamp 1714281807
transform 1 0 2472 0 1 1170
box -8 -3 16 105
use FILL  FILL_2489
timestamp 1714281807
transform 1 0 2464 0 1 1170
box -8 -3 16 105
use FILL  FILL_2490
timestamp 1714281807
transform 1 0 2456 0 1 1170
box -8 -3 16 105
use FILL  FILL_2491
timestamp 1714281807
transform 1 0 2416 0 1 1170
box -8 -3 16 105
use FILL  FILL_2492
timestamp 1714281807
transform 1 0 2352 0 1 1170
box -8 -3 16 105
use FILL  FILL_2493
timestamp 1714281807
transform 1 0 2344 0 1 1170
box -8 -3 16 105
use FILL  FILL_2494
timestamp 1714281807
transform 1 0 2336 0 1 1170
box -8 -3 16 105
use FILL  FILL_2495
timestamp 1714281807
transform 1 0 2328 0 1 1170
box -8 -3 16 105
use FILL  FILL_2496
timestamp 1714281807
transform 1 0 2320 0 1 1170
box -8 -3 16 105
use FILL  FILL_2497
timestamp 1714281807
transform 1 0 2272 0 1 1170
box -8 -3 16 105
use FILL  FILL_2498
timestamp 1714281807
transform 1 0 2264 0 1 1170
box -8 -3 16 105
use FILL  FILL_2499
timestamp 1714281807
transform 1 0 2256 0 1 1170
box -8 -3 16 105
use FILL  FILL_2500
timestamp 1714281807
transform 1 0 2248 0 1 1170
box -8 -3 16 105
use FILL  FILL_2501
timestamp 1714281807
transform 1 0 2240 0 1 1170
box -8 -3 16 105
use FILL  FILL_2502
timestamp 1714281807
transform 1 0 2232 0 1 1170
box -8 -3 16 105
use FILL  FILL_2503
timestamp 1714281807
transform 1 0 2224 0 1 1170
box -8 -3 16 105
use FILL  FILL_2504
timestamp 1714281807
transform 1 0 2184 0 1 1170
box -8 -3 16 105
use FILL  FILL_2505
timestamp 1714281807
transform 1 0 2176 0 1 1170
box -8 -3 16 105
use FILL  FILL_2506
timestamp 1714281807
transform 1 0 2168 0 1 1170
box -8 -3 16 105
use FILL  FILL_2507
timestamp 1714281807
transform 1 0 2160 0 1 1170
box -8 -3 16 105
use FILL  FILL_2508
timestamp 1714281807
transform 1 0 2056 0 1 1170
box -8 -3 16 105
use FILL  FILL_2509
timestamp 1714281807
transform 1 0 2048 0 1 1170
box -8 -3 16 105
use FILL  FILL_2510
timestamp 1714281807
transform 1 0 2040 0 1 1170
box -8 -3 16 105
use FILL  FILL_2511
timestamp 1714281807
transform 1 0 2032 0 1 1170
box -8 -3 16 105
use FILL  FILL_2512
timestamp 1714281807
transform 1 0 2024 0 1 1170
box -8 -3 16 105
use FILL  FILL_2513
timestamp 1714281807
transform 1 0 2016 0 1 1170
box -8 -3 16 105
use FILL  FILL_2514
timestamp 1714281807
transform 1 0 1976 0 1 1170
box -8 -3 16 105
use FILL  FILL_2515
timestamp 1714281807
transform 1 0 1968 0 1 1170
box -8 -3 16 105
use FILL  FILL_2516
timestamp 1714281807
transform 1 0 1960 0 1 1170
box -8 -3 16 105
use FILL  FILL_2517
timestamp 1714281807
transform 1 0 1952 0 1 1170
box -8 -3 16 105
use FILL  FILL_2518
timestamp 1714281807
transform 1 0 1944 0 1 1170
box -8 -3 16 105
use FILL  FILL_2519
timestamp 1714281807
transform 1 0 1920 0 1 1170
box -8 -3 16 105
use FILL  FILL_2520
timestamp 1714281807
transform 1 0 1912 0 1 1170
box -8 -3 16 105
use FILL  FILL_2521
timestamp 1714281807
transform 1 0 1904 0 1 1170
box -8 -3 16 105
use FILL  FILL_2522
timestamp 1714281807
transform 1 0 1896 0 1 1170
box -8 -3 16 105
use FILL  FILL_2523
timestamp 1714281807
transform 1 0 1888 0 1 1170
box -8 -3 16 105
use FILL  FILL_2524
timestamp 1714281807
transform 1 0 1880 0 1 1170
box -8 -3 16 105
use FILL  FILL_2525
timestamp 1714281807
transform 1 0 1872 0 1 1170
box -8 -3 16 105
use FILL  FILL_2526
timestamp 1714281807
transform 1 0 1864 0 1 1170
box -8 -3 16 105
use FILL  FILL_2527
timestamp 1714281807
transform 1 0 1816 0 1 1170
box -8 -3 16 105
use FILL  FILL_2528
timestamp 1714281807
transform 1 0 1808 0 1 1170
box -8 -3 16 105
use FILL  FILL_2529
timestamp 1714281807
transform 1 0 1800 0 1 1170
box -8 -3 16 105
use FILL  FILL_2530
timestamp 1714281807
transform 1 0 1792 0 1 1170
box -8 -3 16 105
use FILL  FILL_2531
timestamp 1714281807
transform 1 0 1784 0 1 1170
box -8 -3 16 105
use FILL  FILL_2532
timestamp 1714281807
transform 1 0 1776 0 1 1170
box -8 -3 16 105
use FILL  FILL_2533
timestamp 1714281807
transform 1 0 1736 0 1 1170
box -8 -3 16 105
use FILL  FILL_2534
timestamp 1714281807
transform 1 0 1728 0 1 1170
box -8 -3 16 105
use FILL  FILL_2535
timestamp 1714281807
transform 1 0 1720 0 1 1170
box -8 -3 16 105
use FILL  FILL_2536
timestamp 1714281807
transform 1 0 1680 0 1 1170
box -8 -3 16 105
use FILL  FILL_2537
timestamp 1714281807
transform 1 0 1672 0 1 1170
box -8 -3 16 105
use FILL  FILL_2538
timestamp 1714281807
transform 1 0 1664 0 1 1170
box -8 -3 16 105
use FILL  FILL_2539
timestamp 1714281807
transform 1 0 1656 0 1 1170
box -8 -3 16 105
use FILL  FILL_2540
timestamp 1714281807
transform 1 0 1648 0 1 1170
box -8 -3 16 105
use FILL  FILL_2541
timestamp 1714281807
transform 1 0 1616 0 1 1170
box -8 -3 16 105
use FILL  FILL_2542
timestamp 1714281807
transform 1 0 1608 0 1 1170
box -8 -3 16 105
use FILL  FILL_2543
timestamp 1714281807
transform 1 0 1504 0 1 1170
box -8 -3 16 105
use FILL  FILL_2544
timestamp 1714281807
transform 1 0 1496 0 1 1170
box -8 -3 16 105
use FILL  FILL_2545
timestamp 1714281807
transform 1 0 1488 0 1 1170
box -8 -3 16 105
use FILL  FILL_2546
timestamp 1714281807
transform 1 0 1480 0 1 1170
box -8 -3 16 105
use FILL  FILL_2547
timestamp 1714281807
transform 1 0 1432 0 1 1170
box -8 -3 16 105
use FILL  FILL_2548
timestamp 1714281807
transform 1 0 1424 0 1 1170
box -8 -3 16 105
use FILL  FILL_2549
timestamp 1714281807
transform 1 0 1416 0 1 1170
box -8 -3 16 105
use FILL  FILL_2550
timestamp 1714281807
transform 1 0 1312 0 1 1170
box -8 -3 16 105
use FILL  FILL_2551
timestamp 1714281807
transform 1 0 1304 0 1 1170
box -8 -3 16 105
use FILL  FILL_2552
timestamp 1714281807
transform 1 0 1296 0 1 1170
box -8 -3 16 105
use FILL  FILL_2553
timestamp 1714281807
transform 1 0 1264 0 1 1170
box -8 -3 16 105
use FILL  FILL_2554
timestamp 1714281807
transform 1 0 1256 0 1 1170
box -8 -3 16 105
use FILL  FILL_2555
timestamp 1714281807
transform 1 0 1176 0 1 1170
box -8 -3 16 105
use FILL  FILL_2556
timestamp 1714281807
transform 1 0 1152 0 1 1170
box -8 -3 16 105
use FILL  FILL_2557
timestamp 1714281807
transform 1 0 1144 0 1 1170
box -8 -3 16 105
use FILL  FILL_2558
timestamp 1714281807
transform 1 0 1136 0 1 1170
box -8 -3 16 105
use FILL  FILL_2559
timestamp 1714281807
transform 1 0 1128 0 1 1170
box -8 -3 16 105
use FILL  FILL_2560
timestamp 1714281807
transform 1 0 1120 0 1 1170
box -8 -3 16 105
use FILL  FILL_2561
timestamp 1714281807
transform 1 0 1088 0 1 1170
box -8 -3 16 105
use FILL  FILL_2562
timestamp 1714281807
transform 1 0 1032 0 1 1170
box -8 -3 16 105
use FILL  FILL_2563
timestamp 1714281807
transform 1 0 1024 0 1 1170
box -8 -3 16 105
use FILL  FILL_2564
timestamp 1714281807
transform 1 0 1016 0 1 1170
box -8 -3 16 105
use FILL  FILL_2565
timestamp 1714281807
transform 1 0 1008 0 1 1170
box -8 -3 16 105
use FILL  FILL_2566
timestamp 1714281807
transform 1 0 976 0 1 1170
box -8 -3 16 105
use FILL  FILL_2567
timestamp 1714281807
transform 1 0 968 0 1 1170
box -8 -3 16 105
use FILL  FILL_2568
timestamp 1714281807
transform 1 0 928 0 1 1170
box -8 -3 16 105
use FILL  FILL_2569
timestamp 1714281807
transform 1 0 920 0 1 1170
box -8 -3 16 105
use FILL  FILL_2570
timestamp 1714281807
transform 1 0 912 0 1 1170
box -8 -3 16 105
use FILL  FILL_2571
timestamp 1714281807
transform 1 0 904 0 1 1170
box -8 -3 16 105
use FILL  FILL_2572
timestamp 1714281807
transform 1 0 896 0 1 1170
box -8 -3 16 105
use FILL  FILL_2573
timestamp 1714281807
transform 1 0 848 0 1 1170
box -8 -3 16 105
use FILL  FILL_2574
timestamp 1714281807
transform 1 0 840 0 1 1170
box -8 -3 16 105
use FILL  FILL_2575
timestamp 1714281807
transform 1 0 832 0 1 1170
box -8 -3 16 105
use FILL  FILL_2576
timestamp 1714281807
transform 1 0 728 0 1 1170
box -8 -3 16 105
use FILL  FILL_2577
timestamp 1714281807
transform 1 0 720 0 1 1170
box -8 -3 16 105
use FILL  FILL_2578
timestamp 1714281807
transform 1 0 712 0 1 1170
box -8 -3 16 105
use FILL  FILL_2579
timestamp 1714281807
transform 1 0 664 0 1 1170
box -8 -3 16 105
use FILL  FILL_2580
timestamp 1714281807
transform 1 0 656 0 1 1170
box -8 -3 16 105
use FILL  FILL_2581
timestamp 1714281807
transform 1 0 648 0 1 1170
box -8 -3 16 105
use FILL  FILL_2582
timestamp 1714281807
transform 1 0 640 0 1 1170
box -8 -3 16 105
use FILL  FILL_2583
timestamp 1714281807
transform 1 0 632 0 1 1170
box -8 -3 16 105
use FILL  FILL_2584
timestamp 1714281807
transform 1 0 624 0 1 1170
box -8 -3 16 105
use FILL  FILL_2585
timestamp 1714281807
transform 1 0 576 0 1 1170
box -8 -3 16 105
use FILL  FILL_2586
timestamp 1714281807
transform 1 0 568 0 1 1170
box -8 -3 16 105
use FILL  FILL_2587
timestamp 1714281807
transform 1 0 560 0 1 1170
box -8 -3 16 105
use FILL  FILL_2588
timestamp 1714281807
transform 1 0 552 0 1 1170
box -8 -3 16 105
use FILL  FILL_2589
timestamp 1714281807
transform 1 0 544 0 1 1170
box -8 -3 16 105
use FILL  FILL_2590
timestamp 1714281807
transform 1 0 496 0 1 1170
box -8 -3 16 105
use FILL  FILL_2591
timestamp 1714281807
transform 1 0 488 0 1 1170
box -8 -3 16 105
use FILL  FILL_2592
timestamp 1714281807
transform 1 0 480 0 1 1170
box -8 -3 16 105
use FILL  FILL_2593
timestamp 1714281807
transform 1 0 472 0 1 1170
box -8 -3 16 105
use FILL  FILL_2594
timestamp 1714281807
transform 1 0 424 0 1 1170
box -8 -3 16 105
use FILL  FILL_2595
timestamp 1714281807
transform 1 0 416 0 1 1170
box -8 -3 16 105
use FILL  FILL_2596
timestamp 1714281807
transform 1 0 408 0 1 1170
box -8 -3 16 105
use FILL  FILL_2597
timestamp 1714281807
transform 1 0 304 0 1 1170
box -8 -3 16 105
use FILL  FILL_2598
timestamp 1714281807
transform 1 0 296 0 1 1170
box -8 -3 16 105
use FILL  FILL_2599
timestamp 1714281807
transform 1 0 256 0 1 1170
box -8 -3 16 105
use FILL  FILL_2600
timestamp 1714281807
transform 1 0 248 0 1 1170
box -8 -3 16 105
use FILL  FILL_2601
timestamp 1714281807
transform 1 0 216 0 1 1170
box -8 -3 16 105
use FILL  FILL_2602
timestamp 1714281807
transform 1 0 208 0 1 1170
box -8 -3 16 105
use FILL  FILL_2603
timestamp 1714281807
transform 1 0 200 0 1 1170
box -8 -3 16 105
use FILL  FILL_2604
timestamp 1714281807
transform 1 0 192 0 1 1170
box -8 -3 16 105
use FILL  FILL_2605
timestamp 1714281807
transform 1 0 88 0 1 1170
box -8 -3 16 105
use FILL  FILL_2606
timestamp 1714281807
transform 1 0 80 0 1 1170
box -8 -3 16 105
use FILL  FILL_2607
timestamp 1714281807
transform 1 0 72 0 1 1170
box -8 -3 16 105
use FILL  FILL_2608
timestamp 1714281807
transform 1 0 3000 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2609
timestamp 1714281807
transform 1 0 2992 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2610
timestamp 1714281807
transform 1 0 2984 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2611
timestamp 1714281807
transform 1 0 2976 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2612
timestamp 1714281807
transform 1 0 2968 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2613
timestamp 1714281807
transform 1 0 2960 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2614
timestamp 1714281807
transform 1 0 2952 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2615
timestamp 1714281807
transform 1 0 2944 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2616
timestamp 1714281807
transform 1 0 2936 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2617
timestamp 1714281807
transform 1 0 2928 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2618
timestamp 1714281807
transform 1 0 2920 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2619
timestamp 1714281807
transform 1 0 2912 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2620
timestamp 1714281807
transform 1 0 2904 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2621
timestamp 1714281807
transform 1 0 2872 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2622
timestamp 1714281807
transform 1 0 2864 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2623
timestamp 1714281807
transform 1 0 2856 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2624
timestamp 1714281807
transform 1 0 2824 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2625
timestamp 1714281807
transform 1 0 2816 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2626
timestamp 1714281807
transform 1 0 2712 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2627
timestamp 1714281807
transform 1 0 2704 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2628
timestamp 1714281807
transform 1 0 2368 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2629
timestamp 1714281807
transform 1 0 2328 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2630
timestamp 1714281807
transform 1 0 2320 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2631
timestamp 1714281807
transform 1 0 2272 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2632
timestamp 1714281807
transform 1 0 2264 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2633
timestamp 1714281807
transform 1 0 2256 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2634
timestamp 1714281807
transform 1 0 2248 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2635
timestamp 1714281807
transform 1 0 2240 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2636
timestamp 1714281807
transform 1 0 2232 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2637
timestamp 1714281807
transform 1 0 2184 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2638
timestamp 1714281807
transform 1 0 2176 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2639
timestamp 1714281807
transform 1 0 2168 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2640
timestamp 1714281807
transform 1 0 2128 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2641
timestamp 1714281807
transform 1 0 2120 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2642
timestamp 1714281807
transform 1 0 2016 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2643
timestamp 1714281807
transform 1 0 1984 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2644
timestamp 1714281807
transform 1 0 1976 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2645
timestamp 1714281807
transform 1 0 1872 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2646
timestamp 1714281807
transform 1 0 1864 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2647
timestamp 1714281807
transform 1 0 1856 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2648
timestamp 1714281807
transform 1 0 1816 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2649
timestamp 1714281807
transform 1 0 1752 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2650
timestamp 1714281807
transform 1 0 1744 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2651
timestamp 1714281807
transform 1 0 1736 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2652
timestamp 1714281807
transform 1 0 1728 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2653
timestamp 1714281807
transform 1 0 1680 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2654
timestamp 1714281807
transform 1 0 1672 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2655
timestamp 1714281807
transform 1 0 1664 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2656
timestamp 1714281807
transform 1 0 1656 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2657
timestamp 1714281807
transform 1 0 1648 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2658
timestamp 1714281807
transform 1 0 1640 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2659
timestamp 1714281807
transform 1 0 1600 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2660
timestamp 1714281807
transform 1 0 1592 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2661
timestamp 1714281807
transform 1 0 1584 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2662
timestamp 1714281807
transform 1 0 1576 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2663
timestamp 1714281807
transform 1 0 1568 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2664
timestamp 1714281807
transform 1 0 1536 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2665
timestamp 1714281807
transform 1 0 1528 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2666
timestamp 1714281807
transform 1 0 1520 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2667
timestamp 1714281807
transform 1 0 1512 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2668
timestamp 1714281807
transform 1 0 1504 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2669
timestamp 1714281807
transform 1 0 1496 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2670
timestamp 1714281807
transform 1 0 1456 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2671
timestamp 1714281807
transform 1 0 1448 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2672
timestamp 1714281807
transform 1 0 1440 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2673
timestamp 1714281807
transform 1 0 1416 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2674
timestamp 1714281807
transform 1 0 1408 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2675
timestamp 1714281807
transform 1 0 1344 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2676
timestamp 1714281807
transform 1 0 1336 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2677
timestamp 1714281807
transform 1 0 1328 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2678
timestamp 1714281807
transform 1 0 1320 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2679
timestamp 1714281807
transform 1 0 1312 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2680
timestamp 1714281807
transform 1 0 1280 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2681
timestamp 1714281807
transform 1 0 1272 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2682
timestamp 1714281807
transform 1 0 1264 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2683
timestamp 1714281807
transform 1 0 1256 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2684
timestamp 1714281807
transform 1 0 1232 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2685
timestamp 1714281807
transform 1 0 1224 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2686
timestamp 1714281807
transform 1 0 1216 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2687
timestamp 1714281807
transform 1 0 1208 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2688
timestamp 1714281807
transform 1 0 1176 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2689
timestamp 1714281807
transform 1 0 1168 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2690
timestamp 1714281807
transform 1 0 1160 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2691
timestamp 1714281807
transform 1 0 1152 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2692
timestamp 1714281807
transform 1 0 1144 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2693
timestamp 1714281807
transform 1 0 1136 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2694
timestamp 1714281807
transform 1 0 1104 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2695
timestamp 1714281807
transform 1 0 1096 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2696
timestamp 1714281807
transform 1 0 1088 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2697
timestamp 1714281807
transform 1 0 1080 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2698
timestamp 1714281807
transform 1 0 1056 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2699
timestamp 1714281807
transform 1 0 1048 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2700
timestamp 1714281807
transform 1 0 1040 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2701
timestamp 1714281807
transform 1 0 992 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2702
timestamp 1714281807
transform 1 0 984 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2703
timestamp 1714281807
transform 1 0 976 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2704
timestamp 1714281807
transform 1 0 936 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2705
timestamp 1714281807
transform 1 0 928 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2706
timestamp 1714281807
transform 1 0 920 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2707
timestamp 1714281807
transform 1 0 912 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2708
timestamp 1714281807
transform 1 0 904 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2709
timestamp 1714281807
transform 1 0 896 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2710
timestamp 1714281807
transform 1 0 848 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2711
timestamp 1714281807
transform 1 0 840 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2712
timestamp 1714281807
transform 1 0 832 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2713
timestamp 1714281807
transform 1 0 824 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2714
timestamp 1714281807
transform 1 0 816 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2715
timestamp 1714281807
transform 1 0 784 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2716
timestamp 1714281807
transform 1 0 776 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2717
timestamp 1714281807
transform 1 0 768 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2718
timestamp 1714281807
transform 1 0 760 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2719
timestamp 1714281807
transform 1 0 728 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2720
timestamp 1714281807
transform 1 0 720 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2721
timestamp 1714281807
transform 1 0 712 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2722
timestamp 1714281807
transform 1 0 704 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2723
timestamp 1714281807
transform 1 0 664 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2724
timestamp 1714281807
transform 1 0 656 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2725
timestamp 1714281807
transform 1 0 648 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2726
timestamp 1714281807
transform 1 0 640 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2727
timestamp 1714281807
transform 1 0 608 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2728
timestamp 1714281807
transform 1 0 600 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2729
timestamp 1714281807
transform 1 0 592 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2730
timestamp 1714281807
transform 1 0 584 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2731
timestamp 1714281807
transform 1 0 576 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2732
timestamp 1714281807
transform 1 0 568 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2733
timestamp 1714281807
transform 1 0 520 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2734
timestamp 1714281807
transform 1 0 512 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2735
timestamp 1714281807
transform 1 0 504 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2736
timestamp 1714281807
transform 1 0 496 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2737
timestamp 1714281807
transform 1 0 488 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2738
timestamp 1714281807
transform 1 0 464 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2739
timestamp 1714281807
transform 1 0 456 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2740
timestamp 1714281807
transform 1 0 352 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2741
timestamp 1714281807
transform 1 0 344 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2742
timestamp 1714281807
transform 1 0 336 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2743
timestamp 1714281807
transform 1 0 328 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2744
timestamp 1714281807
transform 1 0 320 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2745
timestamp 1714281807
transform 1 0 312 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2746
timestamp 1714281807
transform 1 0 304 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2747
timestamp 1714281807
transform 1 0 296 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2748
timestamp 1714281807
transform 1 0 288 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2749
timestamp 1714281807
transform 1 0 264 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2750
timestamp 1714281807
transform 1 0 256 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2751
timestamp 1714281807
transform 1 0 248 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2752
timestamp 1714281807
transform 1 0 240 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2753
timestamp 1714281807
transform 1 0 232 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2754
timestamp 1714281807
transform 1 0 224 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2755
timestamp 1714281807
transform 1 0 216 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2756
timestamp 1714281807
transform 1 0 208 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2757
timestamp 1714281807
transform 1 0 200 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2758
timestamp 1714281807
transform 1 0 192 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2759
timestamp 1714281807
transform 1 0 184 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2760
timestamp 1714281807
transform 1 0 176 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2761
timestamp 1714281807
transform 1 0 168 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2762
timestamp 1714281807
transform 1 0 160 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2763
timestamp 1714281807
transform 1 0 152 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2764
timestamp 1714281807
transform 1 0 144 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2765
timestamp 1714281807
transform 1 0 136 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2766
timestamp 1714281807
transform 1 0 128 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2767
timestamp 1714281807
transform 1 0 120 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2768
timestamp 1714281807
transform 1 0 112 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2769
timestamp 1714281807
transform 1 0 104 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2770
timestamp 1714281807
transform 1 0 96 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2771
timestamp 1714281807
transform 1 0 88 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2772
timestamp 1714281807
transform 1 0 80 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2773
timestamp 1714281807
transform 1 0 72 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2774
timestamp 1714281807
transform 1 0 3000 0 1 970
box -8 -3 16 105
use FILL  FILL_2775
timestamp 1714281807
transform 1 0 2992 0 1 970
box -8 -3 16 105
use FILL  FILL_2776
timestamp 1714281807
transform 1 0 2984 0 1 970
box -8 -3 16 105
use FILL  FILL_2777
timestamp 1714281807
transform 1 0 2976 0 1 970
box -8 -3 16 105
use FILL  FILL_2778
timestamp 1714281807
transform 1 0 2968 0 1 970
box -8 -3 16 105
use FILL  FILL_2779
timestamp 1714281807
transform 1 0 2960 0 1 970
box -8 -3 16 105
use FILL  FILL_2780
timestamp 1714281807
transform 1 0 2952 0 1 970
box -8 -3 16 105
use FILL  FILL_2781
timestamp 1714281807
transform 1 0 2944 0 1 970
box -8 -3 16 105
use FILL  FILL_2782
timestamp 1714281807
transform 1 0 2936 0 1 970
box -8 -3 16 105
use FILL  FILL_2783
timestamp 1714281807
transform 1 0 2928 0 1 970
box -8 -3 16 105
use FILL  FILL_2784
timestamp 1714281807
transform 1 0 2920 0 1 970
box -8 -3 16 105
use FILL  FILL_2785
timestamp 1714281807
transform 1 0 2816 0 1 970
box -8 -3 16 105
use FILL  FILL_2786
timestamp 1714281807
transform 1 0 2808 0 1 970
box -8 -3 16 105
use FILL  FILL_2787
timestamp 1714281807
transform 1 0 2800 0 1 970
box -8 -3 16 105
use FILL  FILL_2788
timestamp 1714281807
transform 1 0 2792 0 1 970
box -8 -3 16 105
use FILL  FILL_2789
timestamp 1714281807
transform 1 0 2784 0 1 970
box -8 -3 16 105
use FILL  FILL_2790
timestamp 1714281807
transform 1 0 2776 0 1 970
box -8 -3 16 105
use FILL  FILL_2791
timestamp 1714281807
transform 1 0 2768 0 1 970
box -8 -3 16 105
use FILL  FILL_2792
timestamp 1714281807
transform 1 0 2728 0 1 970
box -8 -3 16 105
use FILL  FILL_2793
timestamp 1714281807
transform 1 0 2720 0 1 970
box -8 -3 16 105
use FILL  FILL_2794
timestamp 1714281807
transform 1 0 2712 0 1 970
box -8 -3 16 105
use FILL  FILL_2795
timestamp 1714281807
transform 1 0 2608 0 1 970
box -8 -3 16 105
use FILL  FILL_2796
timestamp 1714281807
transform 1 0 2600 0 1 970
box -8 -3 16 105
use FILL  FILL_2797
timestamp 1714281807
transform 1 0 2568 0 1 970
box -8 -3 16 105
use FILL  FILL_2798
timestamp 1714281807
transform 1 0 2464 0 1 970
box -8 -3 16 105
use FILL  FILL_2799
timestamp 1714281807
transform 1 0 2456 0 1 970
box -8 -3 16 105
use FILL  FILL_2800
timestamp 1714281807
transform 1 0 2448 0 1 970
box -8 -3 16 105
use FILL  FILL_2801
timestamp 1714281807
transform 1 0 2440 0 1 970
box -8 -3 16 105
use FILL  FILL_2802
timestamp 1714281807
transform 1 0 2408 0 1 970
box -8 -3 16 105
use FILL  FILL_2803
timestamp 1714281807
transform 1 0 2400 0 1 970
box -8 -3 16 105
use FILL  FILL_2804
timestamp 1714281807
transform 1 0 2392 0 1 970
box -8 -3 16 105
use FILL  FILL_2805
timestamp 1714281807
transform 1 0 2368 0 1 970
box -8 -3 16 105
use FILL  FILL_2806
timestamp 1714281807
transform 1 0 2360 0 1 970
box -8 -3 16 105
use FILL  FILL_2807
timestamp 1714281807
transform 1 0 2352 0 1 970
box -8 -3 16 105
use FILL  FILL_2808
timestamp 1714281807
transform 1 0 2344 0 1 970
box -8 -3 16 105
use FILL  FILL_2809
timestamp 1714281807
transform 1 0 2240 0 1 970
box -8 -3 16 105
use FILL  FILL_2810
timestamp 1714281807
transform 1 0 2232 0 1 970
box -8 -3 16 105
use FILL  FILL_2811
timestamp 1714281807
transform 1 0 2208 0 1 970
box -8 -3 16 105
use FILL  FILL_2812
timestamp 1714281807
transform 1 0 2104 0 1 970
box -8 -3 16 105
use FILL  FILL_2813
timestamp 1714281807
transform 1 0 2048 0 1 970
box -8 -3 16 105
use FILL  FILL_2814
timestamp 1714281807
transform 1 0 2040 0 1 970
box -8 -3 16 105
use FILL  FILL_2815
timestamp 1714281807
transform 1 0 2032 0 1 970
box -8 -3 16 105
use FILL  FILL_2816
timestamp 1714281807
transform 1 0 1832 0 1 970
box -8 -3 16 105
use FILL  FILL_2817
timestamp 1714281807
transform 1 0 1808 0 1 970
box -8 -3 16 105
use FILL  FILL_2818
timestamp 1714281807
transform 1 0 1800 0 1 970
box -8 -3 16 105
use FILL  FILL_2819
timestamp 1714281807
transform 1 0 1792 0 1 970
box -8 -3 16 105
use FILL  FILL_2820
timestamp 1714281807
transform 1 0 1760 0 1 970
box -8 -3 16 105
use FILL  FILL_2821
timestamp 1714281807
transform 1 0 1752 0 1 970
box -8 -3 16 105
use FILL  FILL_2822
timestamp 1714281807
transform 1 0 1696 0 1 970
box -8 -3 16 105
use FILL  FILL_2823
timestamp 1714281807
transform 1 0 1688 0 1 970
box -8 -3 16 105
use FILL  FILL_2824
timestamp 1714281807
transform 1 0 1568 0 1 970
box -8 -3 16 105
use FILL  FILL_2825
timestamp 1714281807
transform 1 0 1560 0 1 970
box -8 -3 16 105
use FILL  FILL_2826
timestamp 1714281807
transform 1 0 1520 0 1 970
box -8 -3 16 105
use FILL  FILL_2827
timestamp 1714281807
transform 1 0 1512 0 1 970
box -8 -3 16 105
use FILL  FILL_2828
timestamp 1714281807
transform 1 0 1384 0 1 970
box -8 -3 16 105
use FILL  FILL_2829
timestamp 1714281807
transform 1 0 1264 0 1 970
box -8 -3 16 105
use FILL  FILL_2830
timestamp 1714281807
transform 1 0 1216 0 1 970
box -8 -3 16 105
use FILL  FILL_2831
timestamp 1714281807
transform 1 0 1208 0 1 970
box -8 -3 16 105
use FILL  FILL_2832
timestamp 1714281807
transform 1 0 1200 0 1 970
box -8 -3 16 105
use FILL  FILL_2833
timestamp 1714281807
transform 1 0 1192 0 1 970
box -8 -3 16 105
use FILL  FILL_2834
timestamp 1714281807
transform 1 0 1184 0 1 970
box -8 -3 16 105
use FILL  FILL_2835
timestamp 1714281807
transform 1 0 1144 0 1 970
box -8 -3 16 105
use FILL  FILL_2836
timestamp 1714281807
transform 1 0 1136 0 1 970
box -8 -3 16 105
use FILL  FILL_2837
timestamp 1714281807
transform 1 0 1128 0 1 970
box -8 -3 16 105
use FILL  FILL_2838
timestamp 1714281807
transform 1 0 1120 0 1 970
box -8 -3 16 105
use FILL  FILL_2839
timestamp 1714281807
transform 1 0 1112 0 1 970
box -8 -3 16 105
use FILL  FILL_2840
timestamp 1714281807
transform 1 0 1080 0 1 970
box -8 -3 16 105
use FILL  FILL_2841
timestamp 1714281807
transform 1 0 1072 0 1 970
box -8 -3 16 105
use FILL  FILL_2842
timestamp 1714281807
transform 1 0 1064 0 1 970
box -8 -3 16 105
use FILL  FILL_2843
timestamp 1714281807
transform 1 0 1040 0 1 970
box -8 -3 16 105
use FILL  FILL_2844
timestamp 1714281807
transform 1 0 1032 0 1 970
box -8 -3 16 105
use FILL  FILL_2845
timestamp 1714281807
transform 1 0 1024 0 1 970
box -8 -3 16 105
use FILL  FILL_2846
timestamp 1714281807
transform 1 0 1016 0 1 970
box -8 -3 16 105
use FILL  FILL_2847
timestamp 1714281807
transform 1 0 912 0 1 970
box -8 -3 16 105
use FILL  FILL_2848
timestamp 1714281807
transform 1 0 904 0 1 970
box -8 -3 16 105
use FILL  FILL_2849
timestamp 1714281807
transform 1 0 896 0 1 970
box -8 -3 16 105
use FILL  FILL_2850
timestamp 1714281807
transform 1 0 856 0 1 970
box -8 -3 16 105
use FILL  FILL_2851
timestamp 1714281807
transform 1 0 848 0 1 970
box -8 -3 16 105
use FILL  FILL_2852
timestamp 1714281807
transform 1 0 840 0 1 970
box -8 -3 16 105
use FILL  FILL_2853
timestamp 1714281807
transform 1 0 832 0 1 970
box -8 -3 16 105
use FILL  FILL_2854
timestamp 1714281807
transform 1 0 824 0 1 970
box -8 -3 16 105
use FILL  FILL_2855
timestamp 1714281807
transform 1 0 816 0 1 970
box -8 -3 16 105
use FILL  FILL_2856
timestamp 1714281807
transform 1 0 808 0 1 970
box -8 -3 16 105
use FILL  FILL_2857
timestamp 1714281807
transform 1 0 800 0 1 970
box -8 -3 16 105
use FILL  FILL_2858
timestamp 1714281807
transform 1 0 792 0 1 970
box -8 -3 16 105
use FILL  FILL_2859
timestamp 1714281807
transform 1 0 768 0 1 970
box -8 -3 16 105
use FILL  FILL_2860
timestamp 1714281807
transform 1 0 760 0 1 970
box -8 -3 16 105
use FILL  FILL_2861
timestamp 1714281807
transform 1 0 752 0 1 970
box -8 -3 16 105
use FILL  FILL_2862
timestamp 1714281807
transform 1 0 744 0 1 970
box -8 -3 16 105
use FILL  FILL_2863
timestamp 1714281807
transform 1 0 736 0 1 970
box -8 -3 16 105
use FILL  FILL_2864
timestamp 1714281807
transform 1 0 728 0 1 970
box -8 -3 16 105
use FILL  FILL_2865
timestamp 1714281807
transform 1 0 720 0 1 970
box -8 -3 16 105
use FILL  FILL_2866
timestamp 1714281807
transform 1 0 712 0 1 970
box -8 -3 16 105
use FILL  FILL_2867
timestamp 1714281807
transform 1 0 656 0 1 970
box -8 -3 16 105
use FILL  FILL_2868
timestamp 1714281807
transform 1 0 648 0 1 970
box -8 -3 16 105
use FILL  FILL_2869
timestamp 1714281807
transform 1 0 640 0 1 970
box -8 -3 16 105
use FILL  FILL_2870
timestamp 1714281807
transform 1 0 632 0 1 970
box -8 -3 16 105
use FILL  FILL_2871
timestamp 1714281807
transform 1 0 624 0 1 970
box -8 -3 16 105
use FILL  FILL_2872
timestamp 1714281807
transform 1 0 592 0 1 970
box -8 -3 16 105
use FILL  FILL_2873
timestamp 1714281807
transform 1 0 584 0 1 970
box -8 -3 16 105
use FILL  FILL_2874
timestamp 1714281807
transform 1 0 576 0 1 970
box -8 -3 16 105
use FILL  FILL_2875
timestamp 1714281807
transform 1 0 568 0 1 970
box -8 -3 16 105
use FILL  FILL_2876
timestamp 1714281807
transform 1 0 560 0 1 970
box -8 -3 16 105
use FILL  FILL_2877
timestamp 1714281807
transform 1 0 512 0 1 970
box -8 -3 16 105
use FILL  FILL_2878
timestamp 1714281807
transform 1 0 504 0 1 970
box -8 -3 16 105
use FILL  FILL_2879
timestamp 1714281807
transform 1 0 496 0 1 970
box -8 -3 16 105
use FILL  FILL_2880
timestamp 1714281807
transform 1 0 488 0 1 970
box -8 -3 16 105
use FILL  FILL_2881
timestamp 1714281807
transform 1 0 480 0 1 970
box -8 -3 16 105
use FILL  FILL_2882
timestamp 1714281807
transform 1 0 456 0 1 970
box -8 -3 16 105
use FILL  FILL_2883
timestamp 1714281807
transform 1 0 352 0 1 970
box -8 -3 16 105
use FILL  FILL_2884
timestamp 1714281807
transform 1 0 344 0 1 970
box -8 -3 16 105
use FILL  FILL_2885
timestamp 1714281807
transform 1 0 336 0 1 970
box -8 -3 16 105
use FILL  FILL_2886
timestamp 1714281807
transform 1 0 232 0 1 970
box -8 -3 16 105
use FILL  FILL_2887
timestamp 1714281807
transform 1 0 224 0 1 970
box -8 -3 16 105
use FILL  FILL_2888
timestamp 1714281807
transform 1 0 216 0 1 970
box -8 -3 16 105
use FILL  FILL_2889
timestamp 1714281807
transform 1 0 208 0 1 970
box -8 -3 16 105
use FILL  FILL_2890
timestamp 1714281807
transform 1 0 200 0 1 970
box -8 -3 16 105
use FILL  FILL_2891
timestamp 1714281807
transform 1 0 192 0 1 970
box -8 -3 16 105
use FILL  FILL_2892
timestamp 1714281807
transform 1 0 184 0 1 970
box -8 -3 16 105
use FILL  FILL_2893
timestamp 1714281807
transform 1 0 176 0 1 970
box -8 -3 16 105
use FILL  FILL_2894
timestamp 1714281807
transform 1 0 168 0 1 970
box -8 -3 16 105
use FILL  FILL_2895
timestamp 1714281807
transform 1 0 160 0 1 970
box -8 -3 16 105
use FILL  FILL_2896
timestamp 1714281807
transform 1 0 152 0 1 970
box -8 -3 16 105
use FILL  FILL_2897
timestamp 1714281807
transform 1 0 144 0 1 970
box -8 -3 16 105
use FILL  FILL_2898
timestamp 1714281807
transform 1 0 136 0 1 970
box -8 -3 16 105
use FILL  FILL_2899
timestamp 1714281807
transform 1 0 128 0 1 970
box -8 -3 16 105
use FILL  FILL_2900
timestamp 1714281807
transform 1 0 120 0 1 970
box -8 -3 16 105
use FILL  FILL_2901
timestamp 1714281807
transform 1 0 112 0 1 970
box -8 -3 16 105
use FILL  FILL_2902
timestamp 1714281807
transform 1 0 104 0 1 970
box -8 -3 16 105
use FILL  FILL_2903
timestamp 1714281807
transform 1 0 96 0 1 970
box -8 -3 16 105
use FILL  FILL_2904
timestamp 1714281807
transform 1 0 88 0 1 970
box -8 -3 16 105
use FILL  FILL_2905
timestamp 1714281807
transform 1 0 80 0 1 970
box -8 -3 16 105
use FILL  FILL_2906
timestamp 1714281807
transform 1 0 72 0 1 970
box -8 -3 16 105
use FILL  FILL_2907
timestamp 1714281807
transform 1 0 3000 0 -1 970
box -8 -3 16 105
use FILL  FILL_2908
timestamp 1714281807
transform 1 0 2992 0 -1 970
box -8 -3 16 105
use FILL  FILL_2909
timestamp 1714281807
transform 1 0 2984 0 -1 970
box -8 -3 16 105
use FILL  FILL_2910
timestamp 1714281807
transform 1 0 2976 0 -1 970
box -8 -3 16 105
use FILL  FILL_2911
timestamp 1714281807
transform 1 0 2968 0 -1 970
box -8 -3 16 105
use FILL  FILL_2912
timestamp 1714281807
transform 1 0 2960 0 -1 970
box -8 -3 16 105
use FILL  FILL_2913
timestamp 1714281807
transform 1 0 2952 0 -1 970
box -8 -3 16 105
use FILL  FILL_2914
timestamp 1714281807
transform 1 0 2944 0 -1 970
box -8 -3 16 105
use FILL  FILL_2915
timestamp 1714281807
transform 1 0 2840 0 -1 970
box -8 -3 16 105
use FILL  FILL_2916
timestamp 1714281807
transform 1 0 2832 0 -1 970
box -8 -3 16 105
use FILL  FILL_2917
timestamp 1714281807
transform 1 0 2824 0 -1 970
box -8 -3 16 105
use FILL  FILL_2918
timestamp 1714281807
transform 1 0 2816 0 -1 970
box -8 -3 16 105
use FILL  FILL_2919
timestamp 1714281807
transform 1 0 2784 0 -1 970
box -8 -3 16 105
use FILL  FILL_2920
timestamp 1714281807
transform 1 0 2776 0 -1 970
box -8 -3 16 105
use FILL  FILL_2921
timestamp 1714281807
transform 1 0 2752 0 -1 970
box -8 -3 16 105
use FILL  FILL_2922
timestamp 1714281807
transform 1 0 2744 0 -1 970
box -8 -3 16 105
use FILL  FILL_2923
timestamp 1714281807
transform 1 0 2736 0 -1 970
box -8 -3 16 105
use FILL  FILL_2924
timestamp 1714281807
transform 1 0 2632 0 -1 970
box -8 -3 16 105
use FILL  FILL_2925
timestamp 1714281807
transform 1 0 2624 0 -1 970
box -8 -3 16 105
use FILL  FILL_2926
timestamp 1714281807
transform 1 0 2616 0 -1 970
box -8 -3 16 105
use FILL  FILL_2927
timestamp 1714281807
transform 1 0 2608 0 -1 970
box -8 -3 16 105
use FILL  FILL_2928
timestamp 1714281807
transform 1 0 2600 0 -1 970
box -8 -3 16 105
use FILL  FILL_2929
timestamp 1714281807
transform 1 0 2592 0 -1 970
box -8 -3 16 105
use FILL  FILL_2930
timestamp 1714281807
transform 1 0 2584 0 -1 970
box -8 -3 16 105
use FILL  FILL_2931
timestamp 1714281807
transform 1 0 2576 0 -1 970
box -8 -3 16 105
use FILL  FILL_2932
timestamp 1714281807
transform 1 0 2568 0 -1 970
box -8 -3 16 105
use FILL  FILL_2933
timestamp 1714281807
transform 1 0 2560 0 -1 970
box -8 -3 16 105
use FILL  FILL_2934
timestamp 1714281807
transform 1 0 2552 0 -1 970
box -8 -3 16 105
use FILL  FILL_2935
timestamp 1714281807
transform 1 0 2544 0 -1 970
box -8 -3 16 105
use FILL  FILL_2936
timestamp 1714281807
transform 1 0 2536 0 -1 970
box -8 -3 16 105
use FILL  FILL_2937
timestamp 1714281807
transform 1 0 2528 0 -1 970
box -8 -3 16 105
use FILL  FILL_2938
timestamp 1714281807
transform 1 0 2520 0 -1 970
box -8 -3 16 105
use FILL  FILL_2939
timestamp 1714281807
transform 1 0 2512 0 -1 970
box -8 -3 16 105
use FILL  FILL_2940
timestamp 1714281807
transform 1 0 2504 0 -1 970
box -8 -3 16 105
use FILL  FILL_2941
timestamp 1714281807
transform 1 0 2496 0 -1 970
box -8 -3 16 105
use FILL  FILL_2942
timestamp 1714281807
transform 1 0 2488 0 -1 970
box -8 -3 16 105
use FILL  FILL_2943
timestamp 1714281807
transform 1 0 2432 0 -1 970
box -8 -3 16 105
use FILL  FILL_2944
timestamp 1714281807
transform 1 0 2424 0 -1 970
box -8 -3 16 105
use FILL  FILL_2945
timestamp 1714281807
transform 1 0 2416 0 -1 970
box -8 -3 16 105
use FILL  FILL_2946
timestamp 1714281807
transform 1 0 2408 0 -1 970
box -8 -3 16 105
use FILL  FILL_2947
timestamp 1714281807
transform 1 0 2400 0 -1 970
box -8 -3 16 105
use FILL  FILL_2948
timestamp 1714281807
transform 1 0 2296 0 -1 970
box -8 -3 16 105
use FILL  FILL_2949
timestamp 1714281807
transform 1 0 2288 0 -1 970
box -8 -3 16 105
use FILL  FILL_2950
timestamp 1714281807
transform 1 0 2280 0 -1 970
box -8 -3 16 105
use FILL  FILL_2951
timestamp 1714281807
transform 1 0 2272 0 -1 970
box -8 -3 16 105
use FILL  FILL_2952
timestamp 1714281807
transform 1 0 2264 0 -1 970
box -8 -3 16 105
use FILL  FILL_2953
timestamp 1714281807
transform 1 0 2240 0 -1 970
box -8 -3 16 105
use FILL  FILL_2954
timestamp 1714281807
transform 1 0 2232 0 -1 970
box -8 -3 16 105
use FILL  FILL_2955
timestamp 1714281807
transform 1 0 2224 0 -1 970
box -8 -3 16 105
use FILL  FILL_2956
timestamp 1714281807
transform 1 0 2216 0 -1 970
box -8 -3 16 105
use FILL  FILL_2957
timestamp 1714281807
transform 1 0 2208 0 -1 970
box -8 -3 16 105
use FILL  FILL_2958
timestamp 1714281807
transform 1 0 2200 0 -1 970
box -8 -3 16 105
use FILL  FILL_2959
timestamp 1714281807
transform 1 0 2192 0 -1 970
box -8 -3 16 105
use FILL  FILL_2960
timestamp 1714281807
transform 1 0 2184 0 -1 970
box -8 -3 16 105
use FILL  FILL_2961
timestamp 1714281807
transform 1 0 2176 0 -1 970
box -8 -3 16 105
use FILL  FILL_2962
timestamp 1714281807
transform 1 0 2072 0 -1 970
box -8 -3 16 105
use FILL  FILL_2963
timestamp 1714281807
transform 1 0 2064 0 -1 970
box -8 -3 16 105
use FILL  FILL_2964
timestamp 1714281807
transform 1 0 2056 0 -1 970
box -8 -3 16 105
use FILL  FILL_2965
timestamp 1714281807
transform 1 0 2024 0 -1 970
box -8 -3 16 105
use FILL  FILL_2966
timestamp 1714281807
transform 1 0 2016 0 -1 970
box -8 -3 16 105
use FILL  FILL_2967
timestamp 1714281807
transform 1 0 2008 0 -1 970
box -8 -3 16 105
use FILL  FILL_2968
timestamp 1714281807
transform 1 0 2000 0 -1 970
box -8 -3 16 105
use FILL  FILL_2969
timestamp 1714281807
transform 1 0 1992 0 -1 970
box -8 -3 16 105
use FILL  FILL_2970
timestamp 1714281807
transform 1 0 1952 0 -1 970
box -8 -3 16 105
use FILL  FILL_2971
timestamp 1714281807
transform 1 0 1944 0 -1 970
box -8 -3 16 105
use FILL  FILL_2972
timestamp 1714281807
transform 1 0 1920 0 -1 970
box -8 -3 16 105
use FILL  FILL_2973
timestamp 1714281807
transform 1 0 1912 0 -1 970
box -8 -3 16 105
use FILL  FILL_2974
timestamp 1714281807
transform 1 0 1904 0 -1 970
box -8 -3 16 105
use FILL  FILL_2975
timestamp 1714281807
transform 1 0 1896 0 -1 970
box -8 -3 16 105
use FILL  FILL_2976
timestamp 1714281807
transform 1 0 1888 0 -1 970
box -8 -3 16 105
use FILL  FILL_2977
timestamp 1714281807
transform 1 0 1848 0 -1 970
box -8 -3 16 105
use FILL  FILL_2978
timestamp 1714281807
transform 1 0 1840 0 -1 970
box -8 -3 16 105
use FILL  FILL_2979
timestamp 1714281807
transform 1 0 1832 0 -1 970
box -8 -3 16 105
use FILL  FILL_2980
timestamp 1714281807
transform 1 0 1824 0 -1 970
box -8 -3 16 105
use FILL  FILL_2981
timestamp 1714281807
transform 1 0 1720 0 -1 970
box -8 -3 16 105
use FILL  FILL_2982
timestamp 1714281807
transform 1 0 1712 0 -1 970
box -8 -3 16 105
use FILL  FILL_2983
timestamp 1714281807
transform 1 0 1704 0 -1 970
box -8 -3 16 105
use FILL  FILL_2984
timestamp 1714281807
transform 1 0 1696 0 -1 970
box -8 -3 16 105
use FILL  FILL_2985
timestamp 1714281807
transform 1 0 1664 0 -1 970
box -8 -3 16 105
use FILL  FILL_2986
timestamp 1714281807
transform 1 0 1656 0 -1 970
box -8 -3 16 105
use FILL  FILL_2987
timestamp 1714281807
transform 1 0 1648 0 -1 970
box -8 -3 16 105
use FILL  FILL_2988
timestamp 1714281807
transform 1 0 1584 0 -1 970
box -8 -3 16 105
use FILL  FILL_2989
timestamp 1714281807
transform 1 0 1552 0 -1 970
box -8 -3 16 105
use FILL  FILL_2990
timestamp 1714281807
transform 1 0 1496 0 -1 970
box -8 -3 16 105
use FILL  FILL_2991
timestamp 1714281807
transform 1 0 1488 0 -1 970
box -8 -3 16 105
use FILL  FILL_2992
timestamp 1714281807
transform 1 0 1480 0 -1 970
box -8 -3 16 105
use FILL  FILL_2993
timestamp 1714281807
transform 1 0 1472 0 -1 970
box -8 -3 16 105
use FILL  FILL_2994
timestamp 1714281807
transform 1 0 1432 0 -1 970
box -8 -3 16 105
use FILL  FILL_2995
timestamp 1714281807
transform 1 0 1424 0 -1 970
box -8 -3 16 105
use FILL  FILL_2996
timestamp 1714281807
transform 1 0 1416 0 -1 970
box -8 -3 16 105
use FILL  FILL_2997
timestamp 1714281807
transform 1 0 1408 0 -1 970
box -8 -3 16 105
use FILL  FILL_2998
timestamp 1714281807
transform 1 0 1304 0 -1 970
box -8 -3 16 105
use FILL  FILL_2999
timestamp 1714281807
transform 1 0 1296 0 -1 970
box -8 -3 16 105
use FILL  FILL_3000
timestamp 1714281807
transform 1 0 1288 0 -1 970
box -8 -3 16 105
use FILL  FILL_3001
timestamp 1714281807
transform 1 0 1280 0 -1 970
box -8 -3 16 105
use FILL  FILL_3002
timestamp 1714281807
transform 1 0 1272 0 -1 970
box -8 -3 16 105
use FILL  FILL_3003
timestamp 1714281807
transform 1 0 1264 0 -1 970
box -8 -3 16 105
use FILL  FILL_3004
timestamp 1714281807
transform 1 0 1256 0 -1 970
box -8 -3 16 105
use FILL  FILL_3005
timestamp 1714281807
transform 1 0 1248 0 -1 970
box -8 -3 16 105
use FILL  FILL_3006
timestamp 1714281807
transform 1 0 1240 0 -1 970
box -8 -3 16 105
use FILL  FILL_3007
timestamp 1714281807
transform 1 0 1200 0 -1 970
box -8 -3 16 105
use FILL  FILL_3008
timestamp 1714281807
transform 1 0 1192 0 -1 970
box -8 -3 16 105
use FILL  FILL_3009
timestamp 1714281807
transform 1 0 1184 0 -1 970
box -8 -3 16 105
use FILL  FILL_3010
timestamp 1714281807
transform 1 0 1176 0 -1 970
box -8 -3 16 105
use FILL  FILL_3011
timestamp 1714281807
transform 1 0 1168 0 -1 970
box -8 -3 16 105
use FILL  FILL_3012
timestamp 1714281807
transform 1 0 1160 0 -1 970
box -8 -3 16 105
use FILL  FILL_3013
timestamp 1714281807
transform 1 0 1056 0 -1 970
box -8 -3 16 105
use FILL  FILL_3014
timestamp 1714281807
transform 1 0 1048 0 -1 970
box -8 -3 16 105
use FILL  FILL_3015
timestamp 1714281807
transform 1 0 1040 0 -1 970
box -8 -3 16 105
use FILL  FILL_3016
timestamp 1714281807
transform 1 0 992 0 -1 970
box -8 -3 16 105
use FILL  FILL_3017
timestamp 1714281807
transform 1 0 984 0 -1 970
box -8 -3 16 105
use FILL  FILL_3018
timestamp 1714281807
transform 1 0 976 0 -1 970
box -8 -3 16 105
use FILL  FILL_3019
timestamp 1714281807
transform 1 0 968 0 -1 970
box -8 -3 16 105
use FILL  FILL_3020
timestamp 1714281807
transform 1 0 960 0 -1 970
box -8 -3 16 105
use FILL  FILL_3021
timestamp 1714281807
transform 1 0 920 0 -1 970
box -8 -3 16 105
use FILL  FILL_3022
timestamp 1714281807
transform 1 0 912 0 -1 970
box -8 -3 16 105
use FILL  FILL_3023
timestamp 1714281807
transform 1 0 904 0 -1 970
box -8 -3 16 105
use FILL  FILL_3024
timestamp 1714281807
transform 1 0 896 0 -1 970
box -8 -3 16 105
use FILL  FILL_3025
timestamp 1714281807
transform 1 0 888 0 -1 970
box -8 -3 16 105
use FILL  FILL_3026
timestamp 1714281807
transform 1 0 848 0 -1 970
box -8 -3 16 105
use FILL  FILL_3027
timestamp 1714281807
transform 1 0 840 0 -1 970
box -8 -3 16 105
use FILL  FILL_3028
timestamp 1714281807
transform 1 0 832 0 -1 970
box -8 -3 16 105
use FILL  FILL_3029
timestamp 1714281807
transform 1 0 824 0 -1 970
box -8 -3 16 105
use FILL  FILL_3030
timestamp 1714281807
transform 1 0 792 0 -1 970
box -8 -3 16 105
use FILL  FILL_3031
timestamp 1714281807
transform 1 0 784 0 -1 970
box -8 -3 16 105
use FILL  FILL_3032
timestamp 1714281807
transform 1 0 760 0 -1 970
box -8 -3 16 105
use FILL  FILL_3033
timestamp 1714281807
transform 1 0 752 0 -1 970
box -8 -3 16 105
use FILL  FILL_3034
timestamp 1714281807
transform 1 0 744 0 -1 970
box -8 -3 16 105
use FILL  FILL_3035
timestamp 1714281807
transform 1 0 736 0 -1 970
box -8 -3 16 105
use FILL  FILL_3036
timestamp 1714281807
transform 1 0 728 0 -1 970
box -8 -3 16 105
use FILL  FILL_3037
timestamp 1714281807
transform 1 0 696 0 -1 970
box -8 -3 16 105
use FILL  FILL_3038
timestamp 1714281807
transform 1 0 688 0 -1 970
box -8 -3 16 105
use FILL  FILL_3039
timestamp 1714281807
transform 1 0 680 0 -1 970
box -8 -3 16 105
use FILL  FILL_3040
timestamp 1714281807
transform 1 0 672 0 -1 970
box -8 -3 16 105
use FILL  FILL_3041
timestamp 1714281807
transform 1 0 664 0 -1 970
box -8 -3 16 105
use FILL  FILL_3042
timestamp 1714281807
transform 1 0 640 0 -1 970
box -8 -3 16 105
use FILL  FILL_3043
timestamp 1714281807
transform 1 0 632 0 -1 970
box -8 -3 16 105
use FILL  FILL_3044
timestamp 1714281807
transform 1 0 624 0 -1 970
box -8 -3 16 105
use FILL  FILL_3045
timestamp 1714281807
transform 1 0 592 0 -1 970
box -8 -3 16 105
use FILL  FILL_3046
timestamp 1714281807
transform 1 0 584 0 -1 970
box -8 -3 16 105
use FILL  FILL_3047
timestamp 1714281807
transform 1 0 576 0 -1 970
box -8 -3 16 105
use FILL  FILL_3048
timestamp 1714281807
transform 1 0 568 0 -1 970
box -8 -3 16 105
use FILL  FILL_3049
timestamp 1714281807
transform 1 0 560 0 -1 970
box -8 -3 16 105
use FILL  FILL_3050
timestamp 1714281807
transform 1 0 552 0 -1 970
box -8 -3 16 105
use FILL  FILL_3051
timestamp 1714281807
transform 1 0 528 0 -1 970
box -8 -3 16 105
use FILL  FILL_3052
timestamp 1714281807
transform 1 0 520 0 -1 970
box -8 -3 16 105
use FILL  FILL_3053
timestamp 1714281807
transform 1 0 488 0 -1 970
box -8 -3 16 105
use FILL  FILL_3054
timestamp 1714281807
transform 1 0 480 0 -1 970
box -8 -3 16 105
use FILL  FILL_3055
timestamp 1714281807
transform 1 0 472 0 -1 970
box -8 -3 16 105
use FILL  FILL_3056
timestamp 1714281807
transform 1 0 464 0 -1 970
box -8 -3 16 105
use FILL  FILL_3057
timestamp 1714281807
transform 1 0 456 0 -1 970
box -8 -3 16 105
use FILL  FILL_3058
timestamp 1714281807
transform 1 0 448 0 -1 970
box -8 -3 16 105
use FILL  FILL_3059
timestamp 1714281807
transform 1 0 440 0 -1 970
box -8 -3 16 105
use FILL  FILL_3060
timestamp 1714281807
transform 1 0 432 0 -1 970
box -8 -3 16 105
use FILL  FILL_3061
timestamp 1714281807
transform 1 0 392 0 -1 970
box -8 -3 16 105
use FILL  FILL_3062
timestamp 1714281807
transform 1 0 384 0 -1 970
box -8 -3 16 105
use FILL  FILL_3063
timestamp 1714281807
transform 1 0 376 0 -1 970
box -8 -3 16 105
use FILL  FILL_3064
timestamp 1714281807
transform 1 0 368 0 -1 970
box -8 -3 16 105
use FILL  FILL_3065
timestamp 1714281807
transform 1 0 360 0 -1 970
box -8 -3 16 105
use FILL  FILL_3066
timestamp 1714281807
transform 1 0 352 0 -1 970
box -8 -3 16 105
use FILL  FILL_3067
timestamp 1714281807
transform 1 0 344 0 -1 970
box -8 -3 16 105
use FILL  FILL_3068
timestamp 1714281807
transform 1 0 336 0 -1 970
box -8 -3 16 105
use FILL  FILL_3069
timestamp 1714281807
transform 1 0 312 0 -1 970
box -8 -3 16 105
use FILL  FILL_3070
timestamp 1714281807
transform 1 0 304 0 -1 970
box -8 -3 16 105
use FILL  FILL_3071
timestamp 1714281807
transform 1 0 296 0 -1 970
box -8 -3 16 105
use FILL  FILL_3072
timestamp 1714281807
transform 1 0 288 0 -1 970
box -8 -3 16 105
use FILL  FILL_3073
timestamp 1714281807
transform 1 0 280 0 -1 970
box -8 -3 16 105
use FILL  FILL_3074
timestamp 1714281807
transform 1 0 272 0 -1 970
box -8 -3 16 105
use FILL  FILL_3075
timestamp 1714281807
transform 1 0 264 0 -1 970
box -8 -3 16 105
use FILL  FILL_3076
timestamp 1714281807
transform 1 0 256 0 -1 970
box -8 -3 16 105
use FILL  FILL_3077
timestamp 1714281807
transform 1 0 248 0 -1 970
box -8 -3 16 105
use FILL  FILL_3078
timestamp 1714281807
transform 1 0 240 0 -1 970
box -8 -3 16 105
use FILL  FILL_3079
timestamp 1714281807
transform 1 0 232 0 -1 970
box -8 -3 16 105
use FILL  FILL_3080
timestamp 1714281807
transform 1 0 224 0 -1 970
box -8 -3 16 105
use FILL  FILL_3081
timestamp 1714281807
transform 1 0 216 0 -1 970
box -8 -3 16 105
use FILL  FILL_3082
timestamp 1714281807
transform 1 0 208 0 -1 970
box -8 -3 16 105
use FILL  FILL_3083
timestamp 1714281807
transform 1 0 200 0 -1 970
box -8 -3 16 105
use FILL  FILL_3084
timestamp 1714281807
transform 1 0 192 0 -1 970
box -8 -3 16 105
use FILL  FILL_3085
timestamp 1714281807
transform 1 0 184 0 -1 970
box -8 -3 16 105
use FILL  FILL_3086
timestamp 1714281807
transform 1 0 176 0 -1 970
box -8 -3 16 105
use FILL  FILL_3087
timestamp 1714281807
transform 1 0 168 0 -1 970
box -8 -3 16 105
use FILL  FILL_3088
timestamp 1714281807
transform 1 0 160 0 -1 970
box -8 -3 16 105
use FILL  FILL_3089
timestamp 1714281807
transform 1 0 152 0 -1 970
box -8 -3 16 105
use FILL  FILL_3090
timestamp 1714281807
transform 1 0 144 0 -1 970
box -8 -3 16 105
use FILL  FILL_3091
timestamp 1714281807
transform 1 0 136 0 -1 970
box -8 -3 16 105
use FILL  FILL_3092
timestamp 1714281807
transform 1 0 128 0 -1 970
box -8 -3 16 105
use FILL  FILL_3093
timestamp 1714281807
transform 1 0 120 0 -1 970
box -8 -3 16 105
use FILL  FILL_3094
timestamp 1714281807
transform 1 0 112 0 -1 970
box -8 -3 16 105
use FILL  FILL_3095
timestamp 1714281807
transform 1 0 104 0 -1 970
box -8 -3 16 105
use FILL  FILL_3096
timestamp 1714281807
transform 1 0 96 0 -1 970
box -8 -3 16 105
use FILL  FILL_3097
timestamp 1714281807
transform 1 0 88 0 -1 970
box -8 -3 16 105
use FILL  FILL_3098
timestamp 1714281807
transform 1 0 80 0 -1 970
box -8 -3 16 105
use FILL  FILL_3099
timestamp 1714281807
transform 1 0 72 0 -1 970
box -8 -3 16 105
use FILL  FILL_3100
timestamp 1714281807
transform 1 0 3000 0 1 770
box -8 -3 16 105
use FILL  FILL_3101
timestamp 1714281807
transform 1 0 2992 0 1 770
box -8 -3 16 105
use FILL  FILL_3102
timestamp 1714281807
transform 1 0 2984 0 1 770
box -8 -3 16 105
use FILL  FILL_3103
timestamp 1714281807
transform 1 0 2976 0 1 770
box -8 -3 16 105
use FILL  FILL_3104
timestamp 1714281807
transform 1 0 2968 0 1 770
box -8 -3 16 105
use FILL  FILL_3105
timestamp 1714281807
transform 1 0 2960 0 1 770
box -8 -3 16 105
use FILL  FILL_3106
timestamp 1714281807
transform 1 0 2952 0 1 770
box -8 -3 16 105
use FILL  FILL_3107
timestamp 1714281807
transform 1 0 2848 0 1 770
box -8 -3 16 105
use FILL  FILL_3108
timestamp 1714281807
transform 1 0 2840 0 1 770
box -8 -3 16 105
use FILL  FILL_3109
timestamp 1714281807
transform 1 0 2808 0 1 770
box -8 -3 16 105
use FILL  FILL_3110
timestamp 1714281807
transform 1 0 2800 0 1 770
box -8 -3 16 105
use FILL  FILL_3111
timestamp 1714281807
transform 1 0 2792 0 1 770
box -8 -3 16 105
use FILL  FILL_3112
timestamp 1714281807
transform 1 0 2784 0 1 770
box -8 -3 16 105
use FILL  FILL_3113
timestamp 1714281807
transform 1 0 2776 0 1 770
box -8 -3 16 105
use FILL  FILL_3114
timestamp 1714281807
transform 1 0 2736 0 1 770
box -8 -3 16 105
use FILL  FILL_3115
timestamp 1714281807
transform 1 0 2728 0 1 770
box -8 -3 16 105
use FILL  FILL_3116
timestamp 1714281807
transform 1 0 2720 0 1 770
box -8 -3 16 105
use FILL  FILL_3117
timestamp 1714281807
transform 1 0 2712 0 1 770
box -8 -3 16 105
use FILL  FILL_3118
timestamp 1714281807
transform 1 0 2704 0 1 770
box -8 -3 16 105
use FILL  FILL_3119
timestamp 1714281807
transform 1 0 2664 0 1 770
box -8 -3 16 105
use FILL  FILL_3120
timestamp 1714281807
transform 1 0 2656 0 1 770
box -8 -3 16 105
use FILL  FILL_3121
timestamp 1714281807
transform 1 0 2648 0 1 770
box -8 -3 16 105
use FILL  FILL_3122
timestamp 1714281807
transform 1 0 2640 0 1 770
box -8 -3 16 105
use FILL  FILL_3123
timestamp 1714281807
transform 1 0 2632 0 1 770
box -8 -3 16 105
use FILL  FILL_3124
timestamp 1714281807
transform 1 0 2528 0 1 770
box -8 -3 16 105
use FILL  FILL_3125
timestamp 1714281807
transform 1 0 2520 0 1 770
box -8 -3 16 105
use FILL  FILL_3126
timestamp 1714281807
transform 1 0 2512 0 1 770
box -8 -3 16 105
use FILL  FILL_3127
timestamp 1714281807
transform 1 0 2504 0 1 770
box -8 -3 16 105
use FILL  FILL_3128
timestamp 1714281807
transform 1 0 2472 0 1 770
box -8 -3 16 105
use FILL  FILL_3129
timestamp 1714281807
transform 1 0 2464 0 1 770
box -8 -3 16 105
use FILL  FILL_3130
timestamp 1714281807
transform 1 0 2456 0 1 770
box -8 -3 16 105
use FILL  FILL_3131
timestamp 1714281807
transform 1 0 2448 0 1 770
box -8 -3 16 105
use FILL  FILL_3132
timestamp 1714281807
transform 1 0 2440 0 1 770
box -8 -3 16 105
use FILL  FILL_3133
timestamp 1714281807
transform 1 0 2336 0 1 770
box -8 -3 16 105
use FILL  FILL_3134
timestamp 1714281807
transform 1 0 2328 0 1 770
box -8 -3 16 105
use FILL  FILL_3135
timestamp 1714281807
transform 1 0 2320 0 1 770
box -8 -3 16 105
use FILL  FILL_3136
timestamp 1714281807
transform 1 0 2280 0 1 770
box -8 -3 16 105
use FILL  FILL_3137
timestamp 1714281807
transform 1 0 2272 0 1 770
box -8 -3 16 105
use FILL  FILL_3138
timestamp 1714281807
transform 1 0 2264 0 1 770
box -8 -3 16 105
use FILL  FILL_3139
timestamp 1714281807
transform 1 0 2256 0 1 770
box -8 -3 16 105
use FILL  FILL_3140
timestamp 1714281807
transform 1 0 2224 0 1 770
box -8 -3 16 105
use FILL  FILL_3141
timestamp 1714281807
transform 1 0 2216 0 1 770
box -8 -3 16 105
use FILL  FILL_3142
timestamp 1714281807
transform 1 0 2208 0 1 770
box -8 -3 16 105
use FILL  FILL_3143
timestamp 1714281807
transform 1 0 2104 0 1 770
box -8 -3 16 105
use FILL  FILL_3144
timestamp 1714281807
transform 1 0 2000 0 1 770
box -8 -3 16 105
use FILL  FILL_3145
timestamp 1714281807
transform 1 0 1992 0 1 770
box -8 -3 16 105
use FILL  FILL_3146
timestamp 1714281807
transform 1 0 1984 0 1 770
box -8 -3 16 105
use FILL  FILL_3147
timestamp 1714281807
transform 1 0 1976 0 1 770
box -8 -3 16 105
use FILL  FILL_3148
timestamp 1714281807
transform 1 0 1944 0 1 770
box -8 -3 16 105
use FILL  FILL_3149
timestamp 1714281807
transform 1 0 1936 0 1 770
box -8 -3 16 105
use FILL  FILL_3150
timestamp 1714281807
transform 1 0 1912 0 1 770
box -8 -3 16 105
use FILL  FILL_3151
timestamp 1714281807
transform 1 0 1904 0 1 770
box -8 -3 16 105
use FILL  FILL_3152
timestamp 1714281807
transform 1 0 1896 0 1 770
box -8 -3 16 105
use FILL  FILL_3153
timestamp 1714281807
transform 1 0 1792 0 1 770
box -8 -3 16 105
use FILL  FILL_3154
timestamp 1714281807
transform 1 0 1784 0 1 770
box -8 -3 16 105
use FILL  FILL_3155
timestamp 1714281807
transform 1 0 1744 0 1 770
box -8 -3 16 105
use FILL  FILL_3156
timestamp 1714281807
transform 1 0 1736 0 1 770
box -8 -3 16 105
use FILL  FILL_3157
timestamp 1714281807
transform 1 0 1728 0 1 770
box -8 -3 16 105
use FILL  FILL_3158
timestamp 1714281807
transform 1 0 1720 0 1 770
box -8 -3 16 105
use FILL  FILL_3159
timestamp 1714281807
transform 1 0 1616 0 1 770
box -8 -3 16 105
use FILL  FILL_3160
timestamp 1714281807
transform 1 0 1512 0 1 770
box -8 -3 16 105
use FILL  FILL_3161
timestamp 1714281807
transform 1 0 1504 0 1 770
box -8 -3 16 105
use FILL  FILL_3162
timestamp 1714281807
transform 1 0 1496 0 1 770
box -8 -3 16 105
use FILL  FILL_3163
timestamp 1714281807
transform 1 0 1464 0 1 770
box -8 -3 16 105
use FILL  FILL_3164
timestamp 1714281807
transform 1 0 1456 0 1 770
box -8 -3 16 105
use FILL  FILL_3165
timestamp 1714281807
transform 1 0 1448 0 1 770
box -8 -3 16 105
use FILL  FILL_3166
timestamp 1714281807
transform 1 0 1424 0 1 770
box -8 -3 16 105
use FILL  FILL_3167
timestamp 1714281807
transform 1 0 1416 0 1 770
box -8 -3 16 105
use FILL  FILL_3168
timestamp 1714281807
transform 1 0 1408 0 1 770
box -8 -3 16 105
use FILL  FILL_3169
timestamp 1714281807
transform 1 0 1400 0 1 770
box -8 -3 16 105
use FILL  FILL_3170
timestamp 1714281807
transform 1 0 1368 0 1 770
box -8 -3 16 105
use FILL  FILL_3171
timestamp 1714281807
transform 1 0 1360 0 1 770
box -8 -3 16 105
use FILL  FILL_3172
timestamp 1714281807
transform 1 0 1352 0 1 770
box -8 -3 16 105
use FILL  FILL_3173
timestamp 1714281807
transform 1 0 1344 0 1 770
box -8 -3 16 105
use FILL  FILL_3174
timestamp 1714281807
transform 1 0 1304 0 1 770
box -8 -3 16 105
use FILL  FILL_3175
timestamp 1714281807
transform 1 0 1296 0 1 770
box -8 -3 16 105
use FILL  FILL_3176
timestamp 1714281807
transform 1 0 1232 0 1 770
box -8 -3 16 105
use FILL  FILL_3177
timestamp 1714281807
transform 1 0 1224 0 1 770
box -8 -3 16 105
use FILL  FILL_3178
timestamp 1714281807
transform 1 0 1216 0 1 770
box -8 -3 16 105
use FILL  FILL_3179
timestamp 1714281807
transform 1 0 1168 0 1 770
box -8 -3 16 105
use FILL  FILL_3180
timestamp 1714281807
transform 1 0 1160 0 1 770
box -8 -3 16 105
use FILL  FILL_3181
timestamp 1714281807
transform 1 0 1152 0 1 770
box -8 -3 16 105
use FILL  FILL_3182
timestamp 1714281807
transform 1 0 1144 0 1 770
box -8 -3 16 105
use FILL  FILL_3183
timestamp 1714281807
transform 1 0 1136 0 1 770
box -8 -3 16 105
use FILL  FILL_3184
timestamp 1714281807
transform 1 0 1096 0 1 770
box -8 -3 16 105
use FILL  FILL_3185
timestamp 1714281807
transform 1 0 1088 0 1 770
box -8 -3 16 105
use FILL  FILL_3186
timestamp 1714281807
transform 1 0 1080 0 1 770
box -8 -3 16 105
use FILL  FILL_3187
timestamp 1714281807
transform 1 0 336 0 1 770
box -8 -3 16 105
use FILL  FILL_3188
timestamp 1714281807
transform 1 0 328 0 1 770
box -8 -3 16 105
use FILL  FILL_3189
timestamp 1714281807
transform 1 0 224 0 1 770
box -8 -3 16 105
use FILL  FILL_3190
timestamp 1714281807
transform 1 0 216 0 1 770
box -8 -3 16 105
use FILL  FILL_3191
timestamp 1714281807
transform 1 0 208 0 1 770
box -8 -3 16 105
use FILL  FILL_3192
timestamp 1714281807
transform 1 0 200 0 1 770
box -8 -3 16 105
use FILL  FILL_3193
timestamp 1714281807
transform 1 0 192 0 1 770
box -8 -3 16 105
use FILL  FILL_3194
timestamp 1714281807
transform 1 0 184 0 1 770
box -8 -3 16 105
use FILL  FILL_3195
timestamp 1714281807
transform 1 0 176 0 1 770
box -8 -3 16 105
use FILL  FILL_3196
timestamp 1714281807
transform 1 0 168 0 1 770
box -8 -3 16 105
use FILL  FILL_3197
timestamp 1714281807
transform 1 0 160 0 1 770
box -8 -3 16 105
use FILL  FILL_3198
timestamp 1714281807
transform 1 0 152 0 1 770
box -8 -3 16 105
use FILL  FILL_3199
timestamp 1714281807
transform 1 0 144 0 1 770
box -8 -3 16 105
use FILL  FILL_3200
timestamp 1714281807
transform 1 0 136 0 1 770
box -8 -3 16 105
use FILL  FILL_3201
timestamp 1714281807
transform 1 0 128 0 1 770
box -8 -3 16 105
use FILL  FILL_3202
timestamp 1714281807
transform 1 0 120 0 1 770
box -8 -3 16 105
use FILL  FILL_3203
timestamp 1714281807
transform 1 0 112 0 1 770
box -8 -3 16 105
use FILL  FILL_3204
timestamp 1714281807
transform 1 0 104 0 1 770
box -8 -3 16 105
use FILL  FILL_3205
timestamp 1714281807
transform 1 0 96 0 1 770
box -8 -3 16 105
use FILL  FILL_3206
timestamp 1714281807
transform 1 0 88 0 1 770
box -8 -3 16 105
use FILL  FILL_3207
timestamp 1714281807
transform 1 0 80 0 1 770
box -8 -3 16 105
use FILL  FILL_3208
timestamp 1714281807
transform 1 0 72 0 1 770
box -8 -3 16 105
use FILL  FILL_3209
timestamp 1714281807
transform 1 0 3000 0 -1 770
box -8 -3 16 105
use FILL  FILL_3210
timestamp 1714281807
transform 1 0 2992 0 -1 770
box -8 -3 16 105
use FILL  FILL_3211
timestamp 1714281807
transform 1 0 2984 0 -1 770
box -8 -3 16 105
use FILL  FILL_3212
timestamp 1714281807
transform 1 0 2976 0 -1 770
box -8 -3 16 105
use FILL  FILL_3213
timestamp 1714281807
transform 1 0 2968 0 -1 770
box -8 -3 16 105
use FILL  FILL_3214
timestamp 1714281807
transform 1 0 2960 0 -1 770
box -8 -3 16 105
use FILL  FILL_3215
timestamp 1714281807
transform 1 0 2952 0 -1 770
box -8 -3 16 105
use FILL  FILL_3216
timestamp 1714281807
transform 1 0 2944 0 -1 770
box -8 -3 16 105
use FILL  FILL_3217
timestamp 1714281807
transform 1 0 2936 0 -1 770
box -8 -3 16 105
use FILL  FILL_3218
timestamp 1714281807
transform 1 0 2928 0 -1 770
box -8 -3 16 105
use FILL  FILL_3219
timestamp 1714281807
transform 1 0 2920 0 -1 770
box -8 -3 16 105
use FILL  FILL_3220
timestamp 1714281807
transform 1 0 2912 0 -1 770
box -8 -3 16 105
use FILL  FILL_3221
timestamp 1714281807
transform 1 0 2904 0 -1 770
box -8 -3 16 105
use FILL  FILL_3222
timestamp 1714281807
transform 1 0 2896 0 -1 770
box -8 -3 16 105
use FILL  FILL_3223
timestamp 1714281807
transform 1 0 2888 0 -1 770
box -8 -3 16 105
use FILL  FILL_3224
timestamp 1714281807
transform 1 0 2864 0 -1 770
box -8 -3 16 105
use FILL  FILL_3225
timestamp 1714281807
transform 1 0 2856 0 -1 770
box -8 -3 16 105
use FILL  FILL_3226
timestamp 1714281807
transform 1 0 2560 0 -1 770
box -8 -3 16 105
use FILL  FILL_3227
timestamp 1714281807
transform 1 0 2552 0 -1 770
box -8 -3 16 105
use FILL  FILL_3228
timestamp 1714281807
transform 1 0 2544 0 -1 770
box -8 -3 16 105
use FILL  FILL_3229
timestamp 1714281807
transform 1 0 2512 0 -1 770
box -8 -3 16 105
use FILL  FILL_3230
timestamp 1714281807
transform 1 0 2504 0 -1 770
box -8 -3 16 105
use FILL  FILL_3231
timestamp 1714281807
transform 1 0 2464 0 -1 770
box -8 -3 16 105
use FILL  FILL_3232
timestamp 1714281807
transform 1 0 2456 0 -1 770
box -8 -3 16 105
use FILL  FILL_3233
timestamp 1714281807
transform 1 0 2448 0 -1 770
box -8 -3 16 105
use FILL  FILL_3234
timestamp 1714281807
transform 1 0 2440 0 -1 770
box -8 -3 16 105
use FILL  FILL_3235
timestamp 1714281807
transform 1 0 2336 0 -1 770
box -8 -3 16 105
use FILL  FILL_3236
timestamp 1714281807
transform 1 0 2328 0 -1 770
box -8 -3 16 105
use FILL  FILL_3237
timestamp 1714281807
transform 1 0 2296 0 -1 770
box -8 -3 16 105
use FILL  FILL_3238
timestamp 1714281807
transform 1 0 2288 0 -1 770
box -8 -3 16 105
use FILL  FILL_3239
timestamp 1714281807
transform 1 0 2280 0 -1 770
box -8 -3 16 105
use FILL  FILL_3240
timestamp 1714281807
transform 1 0 2272 0 -1 770
box -8 -3 16 105
use FILL  FILL_3241
timestamp 1714281807
transform 1 0 2168 0 -1 770
box -8 -3 16 105
use FILL  FILL_3242
timestamp 1714281807
transform 1 0 2064 0 -1 770
box -8 -3 16 105
use FILL  FILL_3243
timestamp 1714281807
transform 1 0 2056 0 -1 770
box -8 -3 16 105
use FILL  FILL_3244
timestamp 1714281807
transform 1 0 2024 0 -1 770
box -8 -3 16 105
use FILL  FILL_3245
timestamp 1714281807
transform 1 0 2016 0 -1 770
box -8 -3 16 105
use FILL  FILL_3246
timestamp 1714281807
transform 1 0 2008 0 -1 770
box -8 -3 16 105
use FILL  FILL_3247
timestamp 1714281807
transform 1 0 2000 0 -1 770
box -8 -3 16 105
use FILL  FILL_3248
timestamp 1714281807
transform 1 0 1992 0 -1 770
box -8 -3 16 105
use FILL  FILL_3249
timestamp 1714281807
transform 1 0 1936 0 -1 770
box -8 -3 16 105
use FILL  FILL_3250
timestamp 1714281807
transform 1 0 1928 0 -1 770
box -8 -3 16 105
use FILL  FILL_3251
timestamp 1714281807
transform 1 0 1920 0 -1 770
box -8 -3 16 105
use FILL  FILL_3252
timestamp 1714281807
transform 1 0 1720 0 -1 770
box -8 -3 16 105
use FILL  FILL_3253
timestamp 1714281807
transform 1 0 1696 0 -1 770
box -8 -3 16 105
use FILL  FILL_3254
timestamp 1714281807
transform 1 0 1664 0 -1 770
box -8 -3 16 105
use FILL  FILL_3255
timestamp 1714281807
transform 1 0 1656 0 -1 770
box -8 -3 16 105
use FILL  FILL_3256
timestamp 1714281807
transform 1 0 1456 0 -1 770
box -8 -3 16 105
use FILL  FILL_3257
timestamp 1714281807
transform 1 0 1424 0 -1 770
box -8 -3 16 105
use FILL  FILL_3258
timestamp 1714281807
transform 1 0 1416 0 -1 770
box -8 -3 16 105
use FILL  FILL_3259
timestamp 1714281807
transform 1 0 1408 0 -1 770
box -8 -3 16 105
use FILL  FILL_3260
timestamp 1714281807
transform 1 0 1368 0 -1 770
box -8 -3 16 105
use FILL  FILL_3261
timestamp 1714281807
transform 1 0 1360 0 -1 770
box -8 -3 16 105
use FILL  FILL_3262
timestamp 1714281807
transform 1 0 1336 0 -1 770
box -8 -3 16 105
use FILL  FILL_3263
timestamp 1714281807
transform 1 0 1232 0 -1 770
box -8 -3 16 105
use FILL  FILL_3264
timestamp 1714281807
transform 1 0 1224 0 -1 770
box -8 -3 16 105
use FILL  FILL_3265
timestamp 1714281807
transform 1 0 1216 0 -1 770
box -8 -3 16 105
use FILL  FILL_3266
timestamp 1714281807
transform 1 0 1208 0 -1 770
box -8 -3 16 105
use FILL  FILL_3267
timestamp 1714281807
transform 1 0 1160 0 -1 770
box -8 -3 16 105
use FILL  FILL_3268
timestamp 1714281807
transform 1 0 1152 0 -1 770
box -8 -3 16 105
use FILL  FILL_3269
timestamp 1714281807
transform 1 0 1144 0 -1 770
box -8 -3 16 105
use FILL  FILL_3270
timestamp 1714281807
transform 1 0 1136 0 -1 770
box -8 -3 16 105
use FILL  FILL_3271
timestamp 1714281807
transform 1 0 1128 0 -1 770
box -8 -3 16 105
use FILL  FILL_3272
timestamp 1714281807
transform 1 0 1120 0 -1 770
box -8 -3 16 105
use FILL  FILL_3273
timestamp 1714281807
transform 1 0 1080 0 -1 770
box -8 -3 16 105
use FILL  FILL_3274
timestamp 1714281807
transform 1 0 1072 0 -1 770
box -8 -3 16 105
use FILL  FILL_3275
timestamp 1714281807
transform 1 0 1064 0 -1 770
box -8 -3 16 105
use FILL  FILL_3276
timestamp 1714281807
transform 1 0 1032 0 -1 770
box -8 -3 16 105
use FILL  FILL_3277
timestamp 1714281807
transform 1 0 1024 0 -1 770
box -8 -3 16 105
use FILL  FILL_3278
timestamp 1714281807
transform 1 0 1016 0 -1 770
box -8 -3 16 105
use FILL  FILL_3279
timestamp 1714281807
transform 1 0 1008 0 -1 770
box -8 -3 16 105
use FILL  FILL_3280
timestamp 1714281807
transform 1 0 904 0 -1 770
box -8 -3 16 105
use FILL  FILL_3281
timestamp 1714281807
transform 1 0 896 0 -1 770
box -8 -3 16 105
use FILL  FILL_3282
timestamp 1714281807
transform 1 0 888 0 -1 770
box -8 -3 16 105
use FILL  FILL_3283
timestamp 1714281807
transform 1 0 880 0 -1 770
box -8 -3 16 105
use FILL  FILL_3284
timestamp 1714281807
transform 1 0 840 0 -1 770
box -8 -3 16 105
use FILL  FILL_3285
timestamp 1714281807
transform 1 0 832 0 -1 770
box -8 -3 16 105
use FILL  FILL_3286
timestamp 1714281807
transform 1 0 824 0 -1 770
box -8 -3 16 105
use FILL  FILL_3287
timestamp 1714281807
transform 1 0 816 0 -1 770
box -8 -3 16 105
use FILL  FILL_3288
timestamp 1714281807
transform 1 0 784 0 -1 770
box -8 -3 16 105
use FILL  FILL_3289
timestamp 1714281807
transform 1 0 776 0 -1 770
box -8 -3 16 105
use FILL  FILL_3290
timestamp 1714281807
transform 1 0 768 0 -1 770
box -8 -3 16 105
use FILL  FILL_3291
timestamp 1714281807
transform 1 0 760 0 -1 770
box -8 -3 16 105
use FILL  FILL_3292
timestamp 1714281807
transform 1 0 720 0 -1 770
box -8 -3 16 105
use FILL  FILL_3293
timestamp 1714281807
transform 1 0 712 0 -1 770
box -8 -3 16 105
use FILL  FILL_3294
timestamp 1714281807
transform 1 0 704 0 -1 770
box -8 -3 16 105
use FILL  FILL_3295
timestamp 1714281807
transform 1 0 672 0 -1 770
box -8 -3 16 105
use FILL  FILL_3296
timestamp 1714281807
transform 1 0 664 0 -1 770
box -8 -3 16 105
use FILL  FILL_3297
timestamp 1714281807
transform 1 0 656 0 -1 770
box -8 -3 16 105
use FILL  FILL_3298
timestamp 1714281807
transform 1 0 648 0 -1 770
box -8 -3 16 105
use FILL  FILL_3299
timestamp 1714281807
transform 1 0 640 0 -1 770
box -8 -3 16 105
use FILL  FILL_3300
timestamp 1714281807
transform 1 0 608 0 -1 770
box -8 -3 16 105
use FILL  FILL_3301
timestamp 1714281807
transform 1 0 600 0 -1 770
box -8 -3 16 105
use FILL  FILL_3302
timestamp 1714281807
transform 1 0 592 0 -1 770
box -8 -3 16 105
use FILL  FILL_3303
timestamp 1714281807
transform 1 0 560 0 -1 770
box -8 -3 16 105
use FILL  FILL_3304
timestamp 1714281807
transform 1 0 552 0 -1 770
box -8 -3 16 105
use FILL  FILL_3305
timestamp 1714281807
transform 1 0 544 0 -1 770
box -8 -3 16 105
use FILL  FILL_3306
timestamp 1714281807
transform 1 0 536 0 -1 770
box -8 -3 16 105
use FILL  FILL_3307
timestamp 1714281807
transform 1 0 528 0 -1 770
box -8 -3 16 105
use FILL  FILL_3308
timestamp 1714281807
transform 1 0 520 0 -1 770
box -8 -3 16 105
use FILL  FILL_3309
timestamp 1714281807
transform 1 0 488 0 -1 770
box -8 -3 16 105
use FILL  FILL_3310
timestamp 1714281807
transform 1 0 480 0 -1 770
box -8 -3 16 105
use FILL  FILL_3311
timestamp 1714281807
transform 1 0 472 0 -1 770
box -8 -3 16 105
use FILL  FILL_3312
timestamp 1714281807
transform 1 0 448 0 -1 770
box -8 -3 16 105
use FILL  FILL_3313
timestamp 1714281807
transform 1 0 440 0 -1 770
box -8 -3 16 105
use FILL  FILL_3314
timestamp 1714281807
transform 1 0 432 0 -1 770
box -8 -3 16 105
use FILL  FILL_3315
timestamp 1714281807
transform 1 0 424 0 -1 770
box -8 -3 16 105
use FILL  FILL_3316
timestamp 1714281807
transform 1 0 392 0 -1 770
box -8 -3 16 105
use FILL  FILL_3317
timestamp 1714281807
transform 1 0 384 0 -1 770
box -8 -3 16 105
use FILL  FILL_3318
timestamp 1714281807
transform 1 0 376 0 -1 770
box -8 -3 16 105
use FILL  FILL_3319
timestamp 1714281807
transform 1 0 368 0 -1 770
box -8 -3 16 105
use FILL  FILL_3320
timestamp 1714281807
transform 1 0 328 0 -1 770
box -8 -3 16 105
use FILL  FILL_3321
timestamp 1714281807
transform 1 0 320 0 -1 770
box -8 -3 16 105
use FILL  FILL_3322
timestamp 1714281807
transform 1 0 312 0 -1 770
box -8 -3 16 105
use FILL  FILL_3323
timestamp 1714281807
transform 1 0 304 0 -1 770
box -8 -3 16 105
use FILL  FILL_3324
timestamp 1714281807
transform 1 0 296 0 -1 770
box -8 -3 16 105
use FILL  FILL_3325
timestamp 1714281807
transform 1 0 288 0 -1 770
box -8 -3 16 105
use FILL  FILL_3326
timestamp 1714281807
transform 1 0 240 0 -1 770
box -8 -3 16 105
use FILL  FILL_3327
timestamp 1714281807
transform 1 0 232 0 -1 770
box -8 -3 16 105
use FILL  FILL_3328
timestamp 1714281807
transform 1 0 224 0 -1 770
box -8 -3 16 105
use FILL  FILL_3329
timestamp 1714281807
transform 1 0 216 0 -1 770
box -8 -3 16 105
use FILL  FILL_3330
timestamp 1714281807
transform 1 0 208 0 -1 770
box -8 -3 16 105
use FILL  FILL_3331
timestamp 1714281807
transform 1 0 200 0 -1 770
box -8 -3 16 105
use FILL  FILL_3332
timestamp 1714281807
transform 1 0 192 0 -1 770
box -8 -3 16 105
use FILL  FILL_3333
timestamp 1714281807
transform 1 0 184 0 -1 770
box -8 -3 16 105
use FILL  FILL_3334
timestamp 1714281807
transform 1 0 176 0 -1 770
box -8 -3 16 105
use FILL  FILL_3335
timestamp 1714281807
transform 1 0 168 0 -1 770
box -8 -3 16 105
use FILL  FILL_3336
timestamp 1714281807
transform 1 0 160 0 -1 770
box -8 -3 16 105
use FILL  FILL_3337
timestamp 1714281807
transform 1 0 152 0 -1 770
box -8 -3 16 105
use FILL  FILL_3338
timestamp 1714281807
transform 1 0 144 0 -1 770
box -8 -3 16 105
use FILL  FILL_3339
timestamp 1714281807
transform 1 0 136 0 -1 770
box -8 -3 16 105
use FILL  FILL_3340
timestamp 1714281807
transform 1 0 128 0 -1 770
box -8 -3 16 105
use FILL  FILL_3341
timestamp 1714281807
transform 1 0 120 0 -1 770
box -8 -3 16 105
use FILL  FILL_3342
timestamp 1714281807
transform 1 0 112 0 -1 770
box -8 -3 16 105
use FILL  FILL_3343
timestamp 1714281807
transform 1 0 104 0 -1 770
box -8 -3 16 105
use FILL  FILL_3344
timestamp 1714281807
transform 1 0 96 0 -1 770
box -8 -3 16 105
use FILL  FILL_3345
timestamp 1714281807
transform 1 0 88 0 -1 770
box -8 -3 16 105
use FILL  FILL_3346
timestamp 1714281807
transform 1 0 80 0 -1 770
box -8 -3 16 105
use FILL  FILL_3347
timestamp 1714281807
transform 1 0 72 0 -1 770
box -8 -3 16 105
use FILL  FILL_3348
timestamp 1714281807
transform 1 0 3000 0 1 570
box -8 -3 16 105
use FILL  FILL_3349
timestamp 1714281807
transform 1 0 2992 0 1 570
box -8 -3 16 105
use FILL  FILL_3350
timestamp 1714281807
transform 1 0 2984 0 1 570
box -8 -3 16 105
use FILL  FILL_3351
timestamp 1714281807
transform 1 0 2976 0 1 570
box -8 -3 16 105
use FILL  FILL_3352
timestamp 1714281807
transform 1 0 2968 0 1 570
box -8 -3 16 105
use FILL  FILL_3353
timestamp 1714281807
transform 1 0 2960 0 1 570
box -8 -3 16 105
use FILL  FILL_3354
timestamp 1714281807
transform 1 0 2952 0 1 570
box -8 -3 16 105
use FILL  FILL_3355
timestamp 1714281807
transform 1 0 2944 0 1 570
box -8 -3 16 105
use FILL  FILL_3356
timestamp 1714281807
transform 1 0 2936 0 1 570
box -8 -3 16 105
use FILL  FILL_3357
timestamp 1714281807
transform 1 0 2928 0 1 570
box -8 -3 16 105
use FILL  FILL_3358
timestamp 1714281807
transform 1 0 2920 0 1 570
box -8 -3 16 105
use FILL  FILL_3359
timestamp 1714281807
transform 1 0 2912 0 1 570
box -8 -3 16 105
use FILL  FILL_3360
timestamp 1714281807
transform 1 0 2904 0 1 570
box -8 -3 16 105
use FILL  FILL_3361
timestamp 1714281807
transform 1 0 2896 0 1 570
box -8 -3 16 105
use FILL  FILL_3362
timestamp 1714281807
transform 1 0 2888 0 1 570
box -8 -3 16 105
use FILL  FILL_3363
timestamp 1714281807
transform 1 0 2880 0 1 570
box -8 -3 16 105
use FILL  FILL_3364
timestamp 1714281807
transform 1 0 2872 0 1 570
box -8 -3 16 105
use FILL  FILL_3365
timestamp 1714281807
transform 1 0 2768 0 1 570
box -8 -3 16 105
use FILL  FILL_3366
timestamp 1714281807
transform 1 0 2760 0 1 570
box -8 -3 16 105
use FILL  FILL_3367
timestamp 1714281807
transform 1 0 2752 0 1 570
box -8 -3 16 105
use FILL  FILL_3368
timestamp 1714281807
transform 1 0 2744 0 1 570
box -8 -3 16 105
use FILL  FILL_3369
timestamp 1714281807
transform 1 0 2696 0 1 570
box -8 -3 16 105
use FILL  FILL_3370
timestamp 1714281807
transform 1 0 2688 0 1 570
box -8 -3 16 105
use FILL  FILL_3371
timestamp 1714281807
transform 1 0 2680 0 1 570
box -8 -3 16 105
use FILL  FILL_3372
timestamp 1714281807
transform 1 0 2672 0 1 570
box -8 -3 16 105
use FILL  FILL_3373
timestamp 1714281807
transform 1 0 2568 0 1 570
box -8 -3 16 105
use FILL  FILL_3374
timestamp 1714281807
transform 1 0 2560 0 1 570
box -8 -3 16 105
use FILL  FILL_3375
timestamp 1714281807
transform 1 0 2440 0 1 570
box -8 -3 16 105
use FILL  FILL_3376
timestamp 1714281807
transform 1 0 2432 0 1 570
box -8 -3 16 105
use FILL  FILL_3377
timestamp 1714281807
transform 1 0 2392 0 1 570
box -8 -3 16 105
use FILL  FILL_3378
timestamp 1714281807
transform 1 0 2384 0 1 570
box -8 -3 16 105
use FILL  FILL_3379
timestamp 1714281807
transform 1 0 2376 0 1 570
box -8 -3 16 105
use FILL  FILL_3380
timestamp 1714281807
transform 1 0 2368 0 1 570
box -8 -3 16 105
use FILL  FILL_3381
timestamp 1714281807
transform 1 0 2360 0 1 570
box -8 -3 16 105
use FILL  FILL_3382
timestamp 1714281807
transform 1 0 2352 0 1 570
box -8 -3 16 105
use FILL  FILL_3383
timestamp 1714281807
transform 1 0 2344 0 1 570
box -8 -3 16 105
use FILL  FILL_3384
timestamp 1714281807
transform 1 0 2304 0 1 570
box -8 -3 16 105
use FILL  FILL_3385
timestamp 1714281807
transform 1 0 2280 0 1 570
box -8 -3 16 105
use FILL  FILL_3386
timestamp 1714281807
transform 1 0 2272 0 1 570
box -8 -3 16 105
use FILL  FILL_3387
timestamp 1714281807
transform 1 0 2264 0 1 570
box -8 -3 16 105
use FILL  FILL_3388
timestamp 1714281807
transform 1 0 2256 0 1 570
box -8 -3 16 105
use FILL  FILL_3389
timestamp 1714281807
transform 1 0 2152 0 1 570
box -8 -3 16 105
use FILL  FILL_3390
timestamp 1714281807
transform 1 0 2144 0 1 570
box -8 -3 16 105
use FILL  FILL_3391
timestamp 1714281807
transform 1 0 2136 0 1 570
box -8 -3 16 105
use FILL  FILL_3392
timestamp 1714281807
transform 1 0 2128 0 1 570
box -8 -3 16 105
use FILL  FILL_3393
timestamp 1714281807
transform 1 0 2096 0 1 570
box -8 -3 16 105
use FILL  FILL_3394
timestamp 1714281807
transform 1 0 2088 0 1 570
box -8 -3 16 105
use FILL  FILL_3395
timestamp 1714281807
transform 1 0 2080 0 1 570
box -8 -3 16 105
use FILL  FILL_3396
timestamp 1714281807
transform 1 0 2072 0 1 570
box -8 -3 16 105
use FILL  FILL_3397
timestamp 1714281807
transform 1 0 2064 0 1 570
box -8 -3 16 105
use FILL  FILL_3398
timestamp 1714281807
transform 1 0 2056 0 1 570
box -8 -3 16 105
use FILL  FILL_3399
timestamp 1714281807
transform 1 0 2048 0 1 570
box -8 -3 16 105
use FILL  FILL_3400
timestamp 1714281807
transform 1 0 2008 0 1 570
box -8 -3 16 105
use FILL  FILL_3401
timestamp 1714281807
transform 1 0 2000 0 1 570
box -8 -3 16 105
use FILL  FILL_3402
timestamp 1714281807
transform 1 0 1992 0 1 570
box -8 -3 16 105
use FILL  FILL_3403
timestamp 1714281807
transform 1 0 1984 0 1 570
box -8 -3 16 105
use FILL  FILL_3404
timestamp 1714281807
transform 1 0 1880 0 1 570
box -8 -3 16 105
use FILL  FILL_3405
timestamp 1714281807
transform 1 0 1872 0 1 570
box -8 -3 16 105
use FILL  FILL_3406
timestamp 1714281807
transform 1 0 1864 0 1 570
box -8 -3 16 105
use FILL  FILL_3407
timestamp 1714281807
transform 1 0 1832 0 1 570
box -8 -3 16 105
use FILL  FILL_3408
timestamp 1714281807
transform 1 0 1824 0 1 570
box -8 -3 16 105
use FILL  FILL_3409
timestamp 1714281807
transform 1 0 1816 0 1 570
box -8 -3 16 105
use FILL  FILL_3410
timestamp 1714281807
transform 1 0 1808 0 1 570
box -8 -3 16 105
use FILL  FILL_3411
timestamp 1714281807
transform 1 0 1768 0 1 570
box -8 -3 16 105
use FILL  FILL_3412
timestamp 1714281807
transform 1 0 1760 0 1 570
box -8 -3 16 105
use FILL  FILL_3413
timestamp 1714281807
transform 1 0 1752 0 1 570
box -8 -3 16 105
use FILL  FILL_3414
timestamp 1714281807
transform 1 0 1624 0 1 570
box -8 -3 16 105
use FILL  FILL_3415
timestamp 1714281807
transform 1 0 1616 0 1 570
box -8 -3 16 105
use FILL  FILL_3416
timestamp 1714281807
transform 1 0 1608 0 1 570
box -8 -3 16 105
use FILL  FILL_3417
timestamp 1714281807
transform 1 0 1504 0 1 570
box -8 -3 16 105
use FILL  FILL_3418
timestamp 1714281807
transform 1 0 1496 0 1 570
box -8 -3 16 105
use FILL  FILL_3419
timestamp 1714281807
transform 1 0 1488 0 1 570
box -8 -3 16 105
use FILL  FILL_3420
timestamp 1714281807
transform 1 0 1456 0 1 570
box -8 -3 16 105
use FILL  FILL_3421
timestamp 1714281807
transform 1 0 1448 0 1 570
box -8 -3 16 105
use FILL  FILL_3422
timestamp 1714281807
transform 1 0 1440 0 1 570
box -8 -3 16 105
use FILL  FILL_3423
timestamp 1714281807
transform 1 0 1432 0 1 570
box -8 -3 16 105
use FILL  FILL_3424
timestamp 1714281807
transform 1 0 1392 0 1 570
box -8 -3 16 105
use FILL  FILL_3425
timestamp 1714281807
transform 1 0 1384 0 1 570
box -8 -3 16 105
use FILL  FILL_3426
timestamp 1714281807
transform 1 0 1376 0 1 570
box -8 -3 16 105
use FILL  FILL_3427
timestamp 1714281807
transform 1 0 1352 0 1 570
box -8 -3 16 105
use FILL  FILL_3428
timestamp 1714281807
transform 1 0 1344 0 1 570
box -8 -3 16 105
use FILL  FILL_3429
timestamp 1714281807
transform 1 0 1240 0 1 570
box -8 -3 16 105
use FILL  FILL_3430
timestamp 1714281807
transform 1 0 1232 0 1 570
box -8 -3 16 105
use FILL  FILL_3431
timestamp 1714281807
transform 1 0 1224 0 1 570
box -8 -3 16 105
use FILL  FILL_3432
timestamp 1714281807
transform 1 0 1216 0 1 570
box -8 -3 16 105
use FILL  FILL_3433
timestamp 1714281807
transform 1 0 1176 0 1 570
box -8 -3 16 105
use FILL  FILL_3434
timestamp 1714281807
transform 1 0 1168 0 1 570
box -8 -3 16 105
use FILL  FILL_3435
timestamp 1714281807
transform 1 0 1104 0 1 570
box -8 -3 16 105
use FILL  FILL_3436
timestamp 1714281807
transform 1 0 1096 0 1 570
box -8 -3 16 105
use FILL  FILL_3437
timestamp 1714281807
transform 1 0 1072 0 1 570
box -8 -3 16 105
use FILL  FILL_3438
timestamp 1714281807
transform 1 0 1064 0 1 570
box -8 -3 16 105
use FILL  FILL_3439
timestamp 1714281807
transform 1 0 1056 0 1 570
box -8 -3 16 105
use FILL  FILL_3440
timestamp 1714281807
transform 1 0 952 0 1 570
box -8 -3 16 105
use FILL  FILL_3441
timestamp 1714281807
transform 1 0 944 0 1 570
box -8 -3 16 105
use FILL  FILL_3442
timestamp 1714281807
transform 1 0 840 0 1 570
box -8 -3 16 105
use FILL  FILL_3443
timestamp 1714281807
transform 1 0 832 0 1 570
box -8 -3 16 105
use FILL  FILL_3444
timestamp 1714281807
transform 1 0 824 0 1 570
box -8 -3 16 105
use FILL  FILL_3445
timestamp 1714281807
transform 1 0 816 0 1 570
box -8 -3 16 105
use FILL  FILL_3446
timestamp 1714281807
transform 1 0 808 0 1 570
box -8 -3 16 105
use FILL  FILL_3447
timestamp 1714281807
transform 1 0 784 0 1 570
box -8 -3 16 105
use FILL  FILL_3448
timestamp 1714281807
transform 1 0 776 0 1 570
box -8 -3 16 105
use FILL  FILL_3449
timestamp 1714281807
transform 1 0 768 0 1 570
box -8 -3 16 105
use FILL  FILL_3450
timestamp 1714281807
transform 1 0 760 0 1 570
box -8 -3 16 105
use FILL  FILL_3451
timestamp 1714281807
transform 1 0 728 0 1 570
box -8 -3 16 105
use FILL  FILL_3452
timestamp 1714281807
transform 1 0 720 0 1 570
box -8 -3 16 105
use FILL  FILL_3453
timestamp 1714281807
transform 1 0 712 0 1 570
box -8 -3 16 105
use FILL  FILL_3454
timestamp 1714281807
transform 1 0 704 0 1 570
box -8 -3 16 105
use FILL  FILL_3455
timestamp 1714281807
transform 1 0 680 0 1 570
box -8 -3 16 105
use FILL  FILL_3456
timestamp 1714281807
transform 1 0 672 0 1 570
box -8 -3 16 105
use FILL  FILL_3457
timestamp 1714281807
transform 1 0 664 0 1 570
box -8 -3 16 105
use FILL  FILL_3458
timestamp 1714281807
transform 1 0 656 0 1 570
box -8 -3 16 105
use FILL  FILL_3459
timestamp 1714281807
transform 1 0 624 0 1 570
box -8 -3 16 105
use FILL  FILL_3460
timestamp 1714281807
transform 1 0 616 0 1 570
box -8 -3 16 105
use FILL  FILL_3461
timestamp 1714281807
transform 1 0 608 0 1 570
box -8 -3 16 105
use FILL  FILL_3462
timestamp 1714281807
transform 1 0 600 0 1 570
box -8 -3 16 105
use FILL  FILL_3463
timestamp 1714281807
transform 1 0 592 0 1 570
box -8 -3 16 105
use FILL  FILL_3464
timestamp 1714281807
transform 1 0 584 0 1 570
box -8 -3 16 105
use FILL  FILL_3465
timestamp 1714281807
transform 1 0 552 0 1 570
box -8 -3 16 105
use FILL  FILL_3466
timestamp 1714281807
transform 1 0 544 0 1 570
box -8 -3 16 105
use FILL  FILL_3467
timestamp 1714281807
transform 1 0 536 0 1 570
box -8 -3 16 105
use FILL  FILL_3468
timestamp 1714281807
transform 1 0 528 0 1 570
box -8 -3 16 105
use FILL  FILL_3469
timestamp 1714281807
transform 1 0 520 0 1 570
box -8 -3 16 105
use FILL  FILL_3470
timestamp 1714281807
transform 1 0 512 0 1 570
box -8 -3 16 105
use FILL  FILL_3471
timestamp 1714281807
transform 1 0 504 0 1 570
box -8 -3 16 105
use FILL  FILL_3472
timestamp 1714281807
transform 1 0 472 0 1 570
box -8 -3 16 105
use FILL  FILL_3473
timestamp 1714281807
transform 1 0 464 0 1 570
box -8 -3 16 105
use FILL  FILL_3474
timestamp 1714281807
transform 1 0 456 0 1 570
box -8 -3 16 105
use FILL  FILL_3475
timestamp 1714281807
transform 1 0 448 0 1 570
box -8 -3 16 105
use FILL  FILL_3476
timestamp 1714281807
transform 1 0 344 0 1 570
box -8 -3 16 105
use FILL  FILL_3477
timestamp 1714281807
transform 1 0 336 0 1 570
box -8 -3 16 105
use FILL  FILL_3478
timestamp 1714281807
transform 1 0 328 0 1 570
box -8 -3 16 105
use FILL  FILL_3479
timestamp 1714281807
transform 1 0 224 0 1 570
box -8 -3 16 105
use FILL  FILL_3480
timestamp 1714281807
transform 1 0 216 0 1 570
box -8 -3 16 105
use FILL  FILL_3481
timestamp 1714281807
transform 1 0 208 0 1 570
box -8 -3 16 105
use FILL  FILL_3482
timestamp 1714281807
transform 1 0 200 0 1 570
box -8 -3 16 105
use FILL  FILL_3483
timestamp 1714281807
transform 1 0 192 0 1 570
box -8 -3 16 105
use FILL  FILL_3484
timestamp 1714281807
transform 1 0 184 0 1 570
box -8 -3 16 105
use FILL  FILL_3485
timestamp 1714281807
transform 1 0 176 0 1 570
box -8 -3 16 105
use FILL  FILL_3486
timestamp 1714281807
transform 1 0 168 0 1 570
box -8 -3 16 105
use FILL  FILL_3487
timestamp 1714281807
transform 1 0 160 0 1 570
box -8 -3 16 105
use FILL  FILL_3488
timestamp 1714281807
transform 1 0 152 0 1 570
box -8 -3 16 105
use FILL  FILL_3489
timestamp 1714281807
transform 1 0 144 0 1 570
box -8 -3 16 105
use FILL  FILL_3490
timestamp 1714281807
transform 1 0 136 0 1 570
box -8 -3 16 105
use FILL  FILL_3491
timestamp 1714281807
transform 1 0 128 0 1 570
box -8 -3 16 105
use FILL  FILL_3492
timestamp 1714281807
transform 1 0 120 0 1 570
box -8 -3 16 105
use FILL  FILL_3493
timestamp 1714281807
transform 1 0 112 0 1 570
box -8 -3 16 105
use FILL  FILL_3494
timestamp 1714281807
transform 1 0 104 0 1 570
box -8 -3 16 105
use FILL  FILL_3495
timestamp 1714281807
transform 1 0 96 0 1 570
box -8 -3 16 105
use FILL  FILL_3496
timestamp 1714281807
transform 1 0 88 0 1 570
box -8 -3 16 105
use FILL  FILL_3497
timestamp 1714281807
transform 1 0 80 0 1 570
box -8 -3 16 105
use FILL  FILL_3498
timestamp 1714281807
transform 1 0 72 0 1 570
box -8 -3 16 105
use FILL  FILL_3499
timestamp 1714281807
transform 1 0 3000 0 -1 570
box -8 -3 16 105
use FILL  FILL_3500
timestamp 1714281807
transform 1 0 2896 0 -1 570
box -8 -3 16 105
use FILL  FILL_3501
timestamp 1714281807
transform 1 0 2888 0 -1 570
box -8 -3 16 105
use FILL  FILL_3502
timestamp 1714281807
transform 1 0 2864 0 -1 570
box -8 -3 16 105
use FILL  FILL_3503
timestamp 1714281807
transform 1 0 2824 0 -1 570
box -8 -3 16 105
use FILL  FILL_3504
timestamp 1714281807
transform 1 0 2816 0 -1 570
box -8 -3 16 105
use FILL  FILL_3505
timestamp 1714281807
transform 1 0 2808 0 -1 570
box -8 -3 16 105
use FILL  FILL_3506
timestamp 1714281807
transform 1 0 2800 0 -1 570
box -8 -3 16 105
use FILL  FILL_3507
timestamp 1714281807
transform 1 0 2792 0 -1 570
box -8 -3 16 105
use FILL  FILL_3508
timestamp 1714281807
transform 1 0 2784 0 -1 570
box -8 -3 16 105
use FILL  FILL_3509
timestamp 1714281807
transform 1 0 2736 0 -1 570
box -8 -3 16 105
use FILL  FILL_3510
timestamp 1714281807
transform 1 0 2728 0 -1 570
box -8 -3 16 105
use FILL  FILL_3511
timestamp 1714281807
transform 1 0 2720 0 -1 570
box -8 -3 16 105
use FILL  FILL_3512
timestamp 1714281807
transform 1 0 2712 0 -1 570
box -8 -3 16 105
use FILL  FILL_3513
timestamp 1714281807
transform 1 0 2648 0 -1 570
box -8 -3 16 105
use FILL  FILL_3514
timestamp 1714281807
transform 1 0 2640 0 -1 570
box -8 -3 16 105
use FILL  FILL_3515
timestamp 1714281807
transform 1 0 2600 0 -1 570
box -8 -3 16 105
use FILL  FILL_3516
timestamp 1714281807
transform 1 0 2592 0 -1 570
box -8 -3 16 105
use FILL  FILL_3517
timestamp 1714281807
transform 1 0 2584 0 -1 570
box -8 -3 16 105
use FILL  FILL_3518
timestamp 1714281807
transform 1 0 2576 0 -1 570
box -8 -3 16 105
use FILL  FILL_3519
timestamp 1714281807
transform 1 0 2544 0 -1 570
box -8 -3 16 105
use FILL  FILL_3520
timestamp 1714281807
transform 1 0 2536 0 -1 570
box -8 -3 16 105
use FILL  FILL_3521
timestamp 1714281807
transform 1 0 2528 0 -1 570
box -8 -3 16 105
use FILL  FILL_3522
timestamp 1714281807
transform 1 0 2520 0 -1 570
box -8 -3 16 105
use FILL  FILL_3523
timestamp 1714281807
transform 1 0 2512 0 -1 570
box -8 -3 16 105
use FILL  FILL_3524
timestamp 1714281807
transform 1 0 2488 0 -1 570
box -8 -3 16 105
use FILL  FILL_3525
timestamp 1714281807
transform 1 0 2480 0 -1 570
box -8 -3 16 105
use FILL  FILL_3526
timestamp 1714281807
transform 1 0 2472 0 -1 570
box -8 -3 16 105
use FILL  FILL_3527
timestamp 1714281807
transform 1 0 2368 0 -1 570
box -8 -3 16 105
use FILL  FILL_3528
timestamp 1714281807
transform 1 0 2360 0 -1 570
box -8 -3 16 105
use FILL  FILL_3529
timestamp 1714281807
transform 1 0 2256 0 -1 570
box -8 -3 16 105
use FILL  FILL_3530
timestamp 1714281807
transform 1 0 2248 0 -1 570
box -8 -3 16 105
use FILL  FILL_3531
timestamp 1714281807
transform 1 0 2240 0 -1 570
box -8 -3 16 105
use FILL  FILL_3532
timestamp 1714281807
transform 1 0 2232 0 -1 570
box -8 -3 16 105
use FILL  FILL_3533
timestamp 1714281807
transform 1 0 2224 0 -1 570
box -8 -3 16 105
use FILL  FILL_3534
timestamp 1714281807
transform 1 0 2192 0 -1 570
box -8 -3 16 105
use FILL  FILL_3535
timestamp 1714281807
transform 1 0 2184 0 -1 570
box -8 -3 16 105
use FILL  FILL_3536
timestamp 1714281807
transform 1 0 2176 0 -1 570
box -8 -3 16 105
use FILL  FILL_3537
timestamp 1714281807
transform 1 0 2152 0 -1 570
box -8 -3 16 105
use FILL  FILL_3538
timestamp 1714281807
transform 1 0 2144 0 -1 570
box -8 -3 16 105
use FILL  FILL_3539
timestamp 1714281807
transform 1 0 2136 0 -1 570
box -8 -3 16 105
use FILL  FILL_3540
timestamp 1714281807
transform 1 0 2128 0 -1 570
box -8 -3 16 105
use FILL  FILL_3541
timestamp 1714281807
transform 1 0 2120 0 -1 570
box -8 -3 16 105
use FILL  FILL_3542
timestamp 1714281807
transform 1 0 2080 0 -1 570
box -8 -3 16 105
use FILL  FILL_3543
timestamp 1714281807
transform 1 0 2072 0 -1 570
box -8 -3 16 105
use FILL  FILL_3544
timestamp 1714281807
transform 1 0 2064 0 -1 570
box -8 -3 16 105
use FILL  FILL_3545
timestamp 1714281807
transform 1 0 2056 0 -1 570
box -8 -3 16 105
use FILL  FILL_3546
timestamp 1714281807
transform 1 0 2032 0 -1 570
box -8 -3 16 105
use FILL  FILL_3547
timestamp 1714281807
transform 1 0 2024 0 -1 570
box -8 -3 16 105
use FILL  FILL_3548
timestamp 1714281807
transform 1 0 2016 0 -1 570
box -8 -3 16 105
use FILL  FILL_3549
timestamp 1714281807
transform 1 0 1912 0 -1 570
box -8 -3 16 105
use FILL  FILL_3550
timestamp 1714281807
transform 1 0 1904 0 -1 570
box -8 -3 16 105
use FILL  FILL_3551
timestamp 1714281807
transform 1 0 1896 0 -1 570
box -8 -3 16 105
use FILL  FILL_3552
timestamp 1714281807
transform 1 0 1792 0 -1 570
box -8 -3 16 105
use FILL  FILL_3553
timestamp 1714281807
transform 1 0 1784 0 -1 570
box -8 -3 16 105
use FILL  FILL_3554
timestamp 1714281807
transform 1 0 1760 0 -1 570
box -8 -3 16 105
use FILL  FILL_3555
timestamp 1714281807
transform 1 0 1752 0 -1 570
box -8 -3 16 105
use FILL  FILL_3556
timestamp 1714281807
transform 1 0 1744 0 -1 570
box -8 -3 16 105
use FILL  FILL_3557
timestamp 1714281807
transform 1 0 1736 0 -1 570
box -8 -3 16 105
use FILL  FILL_3558
timestamp 1714281807
transform 1 0 1728 0 -1 570
box -8 -3 16 105
use FILL  FILL_3559
timestamp 1714281807
transform 1 0 1720 0 -1 570
box -8 -3 16 105
use FILL  FILL_3560
timestamp 1714281807
transform 1 0 1712 0 -1 570
box -8 -3 16 105
use FILL  FILL_3561
timestamp 1714281807
transform 1 0 1704 0 -1 570
box -8 -3 16 105
use FILL  FILL_3562
timestamp 1714281807
transform 1 0 1664 0 -1 570
box -8 -3 16 105
use FILL  FILL_3563
timestamp 1714281807
transform 1 0 1656 0 -1 570
box -8 -3 16 105
use FILL  FILL_3564
timestamp 1714281807
transform 1 0 1632 0 -1 570
box -8 -3 16 105
use FILL  FILL_3565
timestamp 1714281807
transform 1 0 1624 0 -1 570
box -8 -3 16 105
use FILL  FILL_3566
timestamp 1714281807
transform 1 0 1616 0 -1 570
box -8 -3 16 105
use FILL  FILL_3567
timestamp 1714281807
transform 1 0 1512 0 -1 570
box -8 -3 16 105
use FILL  FILL_3568
timestamp 1714281807
transform 1 0 1504 0 -1 570
box -8 -3 16 105
use FILL  FILL_3569
timestamp 1714281807
transform 1 0 1496 0 -1 570
box -8 -3 16 105
use FILL  FILL_3570
timestamp 1714281807
transform 1 0 1464 0 -1 570
box -8 -3 16 105
use FILL  FILL_3571
timestamp 1714281807
transform 1 0 1456 0 -1 570
box -8 -3 16 105
use FILL  FILL_3572
timestamp 1714281807
transform 1 0 1448 0 -1 570
box -8 -3 16 105
use FILL  FILL_3573
timestamp 1714281807
transform 1 0 1440 0 -1 570
box -8 -3 16 105
use FILL  FILL_3574
timestamp 1714281807
transform 1 0 1432 0 -1 570
box -8 -3 16 105
use FILL  FILL_3575
timestamp 1714281807
transform 1 0 1392 0 -1 570
box -8 -3 16 105
use FILL  FILL_3576
timestamp 1714281807
transform 1 0 1384 0 -1 570
box -8 -3 16 105
use FILL  FILL_3577
timestamp 1714281807
transform 1 0 1360 0 -1 570
box -8 -3 16 105
use FILL  FILL_3578
timestamp 1714281807
transform 1 0 1352 0 -1 570
box -8 -3 16 105
use FILL  FILL_3579
timestamp 1714281807
transform 1 0 1192 0 -1 570
box -8 -3 16 105
use FILL  FILL_3580
timestamp 1714281807
transform 1 0 1184 0 -1 570
box -8 -3 16 105
use FILL  FILL_3581
timestamp 1714281807
transform 1 0 1120 0 -1 570
box -8 -3 16 105
use FILL  FILL_3582
timestamp 1714281807
transform 1 0 1112 0 -1 570
box -8 -3 16 105
use FILL  FILL_3583
timestamp 1714281807
transform 1 0 1104 0 -1 570
box -8 -3 16 105
use FILL  FILL_3584
timestamp 1714281807
transform 1 0 1096 0 -1 570
box -8 -3 16 105
use FILL  FILL_3585
timestamp 1714281807
transform 1 0 1064 0 -1 570
box -8 -3 16 105
use FILL  FILL_3586
timestamp 1714281807
transform 1 0 1056 0 -1 570
box -8 -3 16 105
use FILL  FILL_3587
timestamp 1714281807
transform 1 0 1048 0 -1 570
box -8 -3 16 105
use FILL  FILL_3588
timestamp 1714281807
transform 1 0 944 0 -1 570
box -8 -3 16 105
use FILL  FILL_3589
timestamp 1714281807
transform 1 0 936 0 -1 570
box -8 -3 16 105
use FILL  FILL_3590
timestamp 1714281807
transform 1 0 928 0 -1 570
box -8 -3 16 105
use FILL  FILL_3591
timestamp 1714281807
transform 1 0 920 0 -1 570
box -8 -3 16 105
use FILL  FILL_3592
timestamp 1714281807
transform 1 0 912 0 -1 570
box -8 -3 16 105
use FILL  FILL_3593
timestamp 1714281807
transform 1 0 880 0 -1 570
box -8 -3 16 105
use FILL  FILL_3594
timestamp 1714281807
transform 1 0 872 0 -1 570
box -8 -3 16 105
use FILL  FILL_3595
timestamp 1714281807
transform 1 0 864 0 -1 570
box -8 -3 16 105
use FILL  FILL_3596
timestamp 1714281807
transform 1 0 856 0 -1 570
box -8 -3 16 105
use FILL  FILL_3597
timestamp 1714281807
transform 1 0 752 0 -1 570
box -8 -3 16 105
use FILL  FILL_3598
timestamp 1714281807
transform 1 0 744 0 -1 570
box -8 -3 16 105
use FILL  FILL_3599
timestamp 1714281807
transform 1 0 736 0 -1 570
box -8 -3 16 105
use FILL  FILL_3600
timestamp 1714281807
transform 1 0 728 0 -1 570
box -8 -3 16 105
use FILL  FILL_3601
timestamp 1714281807
transform 1 0 720 0 -1 570
box -8 -3 16 105
use FILL  FILL_3602
timestamp 1714281807
transform 1 0 688 0 -1 570
box -8 -3 16 105
use FILL  FILL_3603
timestamp 1714281807
transform 1 0 680 0 -1 570
box -8 -3 16 105
use FILL  FILL_3604
timestamp 1714281807
transform 1 0 672 0 -1 570
box -8 -3 16 105
use FILL  FILL_3605
timestamp 1714281807
transform 1 0 664 0 -1 570
box -8 -3 16 105
use FILL  FILL_3606
timestamp 1714281807
transform 1 0 656 0 -1 570
box -8 -3 16 105
use FILL  FILL_3607
timestamp 1714281807
transform 1 0 552 0 -1 570
box -8 -3 16 105
use FILL  FILL_3608
timestamp 1714281807
transform 1 0 544 0 -1 570
box -8 -3 16 105
use FILL  FILL_3609
timestamp 1714281807
transform 1 0 536 0 -1 570
box -8 -3 16 105
use FILL  FILL_3610
timestamp 1714281807
transform 1 0 528 0 -1 570
box -8 -3 16 105
use FILL  FILL_3611
timestamp 1714281807
transform 1 0 496 0 -1 570
box -8 -3 16 105
use FILL  FILL_3612
timestamp 1714281807
transform 1 0 488 0 -1 570
box -8 -3 16 105
use FILL  FILL_3613
timestamp 1714281807
transform 1 0 480 0 -1 570
box -8 -3 16 105
use FILL  FILL_3614
timestamp 1714281807
transform 1 0 472 0 -1 570
box -8 -3 16 105
use FILL  FILL_3615
timestamp 1714281807
transform 1 0 464 0 -1 570
box -8 -3 16 105
use FILL  FILL_3616
timestamp 1714281807
transform 1 0 424 0 -1 570
box -8 -3 16 105
use FILL  FILL_3617
timestamp 1714281807
transform 1 0 416 0 -1 570
box -8 -3 16 105
use FILL  FILL_3618
timestamp 1714281807
transform 1 0 408 0 -1 570
box -8 -3 16 105
use FILL  FILL_3619
timestamp 1714281807
transform 1 0 400 0 -1 570
box -8 -3 16 105
use FILL  FILL_3620
timestamp 1714281807
transform 1 0 392 0 -1 570
box -8 -3 16 105
use FILL  FILL_3621
timestamp 1714281807
transform 1 0 288 0 -1 570
box -8 -3 16 105
use FILL  FILL_3622
timestamp 1714281807
transform 1 0 280 0 -1 570
box -8 -3 16 105
use FILL  FILL_3623
timestamp 1714281807
transform 1 0 272 0 -1 570
box -8 -3 16 105
use FILL  FILL_3624
timestamp 1714281807
transform 1 0 264 0 -1 570
box -8 -3 16 105
use FILL  FILL_3625
timestamp 1714281807
transform 1 0 256 0 -1 570
box -8 -3 16 105
use FILL  FILL_3626
timestamp 1714281807
transform 1 0 248 0 -1 570
box -8 -3 16 105
use FILL  FILL_3627
timestamp 1714281807
transform 1 0 240 0 -1 570
box -8 -3 16 105
use FILL  FILL_3628
timestamp 1714281807
transform 1 0 232 0 -1 570
box -8 -3 16 105
use FILL  FILL_3629
timestamp 1714281807
transform 1 0 224 0 -1 570
box -8 -3 16 105
use FILL  FILL_3630
timestamp 1714281807
transform 1 0 216 0 -1 570
box -8 -3 16 105
use FILL  FILL_3631
timestamp 1714281807
transform 1 0 208 0 -1 570
box -8 -3 16 105
use FILL  FILL_3632
timestamp 1714281807
transform 1 0 200 0 -1 570
box -8 -3 16 105
use FILL  FILL_3633
timestamp 1714281807
transform 1 0 192 0 -1 570
box -8 -3 16 105
use FILL  FILL_3634
timestamp 1714281807
transform 1 0 184 0 -1 570
box -8 -3 16 105
use FILL  FILL_3635
timestamp 1714281807
transform 1 0 176 0 -1 570
box -8 -3 16 105
use FILL  FILL_3636
timestamp 1714281807
transform 1 0 168 0 -1 570
box -8 -3 16 105
use FILL  FILL_3637
timestamp 1714281807
transform 1 0 160 0 -1 570
box -8 -3 16 105
use FILL  FILL_3638
timestamp 1714281807
transform 1 0 152 0 -1 570
box -8 -3 16 105
use FILL  FILL_3639
timestamp 1714281807
transform 1 0 144 0 -1 570
box -8 -3 16 105
use FILL  FILL_3640
timestamp 1714281807
transform 1 0 136 0 -1 570
box -8 -3 16 105
use FILL  FILL_3641
timestamp 1714281807
transform 1 0 128 0 -1 570
box -8 -3 16 105
use FILL  FILL_3642
timestamp 1714281807
transform 1 0 120 0 -1 570
box -8 -3 16 105
use FILL  FILL_3643
timestamp 1714281807
transform 1 0 112 0 -1 570
box -8 -3 16 105
use FILL  FILL_3644
timestamp 1714281807
transform 1 0 104 0 -1 570
box -8 -3 16 105
use FILL  FILL_3645
timestamp 1714281807
transform 1 0 96 0 -1 570
box -8 -3 16 105
use FILL  FILL_3646
timestamp 1714281807
transform 1 0 88 0 -1 570
box -8 -3 16 105
use FILL  FILL_3647
timestamp 1714281807
transform 1 0 80 0 -1 570
box -8 -3 16 105
use FILL  FILL_3648
timestamp 1714281807
transform 1 0 72 0 -1 570
box -8 -3 16 105
use FILL  FILL_3649
timestamp 1714281807
transform 1 0 3000 0 1 370
box -8 -3 16 105
use FILL  FILL_3650
timestamp 1714281807
transform 1 0 2992 0 1 370
box -8 -3 16 105
use FILL  FILL_3651
timestamp 1714281807
transform 1 0 2984 0 1 370
box -8 -3 16 105
use FILL  FILL_3652
timestamp 1714281807
transform 1 0 2976 0 1 370
box -8 -3 16 105
use FILL  FILL_3653
timestamp 1714281807
transform 1 0 2968 0 1 370
box -8 -3 16 105
use FILL  FILL_3654
timestamp 1714281807
transform 1 0 2960 0 1 370
box -8 -3 16 105
use FILL  FILL_3655
timestamp 1714281807
transform 1 0 2952 0 1 370
box -8 -3 16 105
use FILL  FILL_3656
timestamp 1714281807
transform 1 0 2944 0 1 370
box -8 -3 16 105
use FILL  FILL_3657
timestamp 1714281807
transform 1 0 2936 0 1 370
box -8 -3 16 105
use FILL  FILL_3658
timestamp 1714281807
transform 1 0 2928 0 1 370
box -8 -3 16 105
use FILL  FILL_3659
timestamp 1714281807
transform 1 0 2864 0 1 370
box -8 -3 16 105
use FILL  FILL_3660
timestamp 1714281807
transform 1 0 2856 0 1 370
box -8 -3 16 105
use FILL  FILL_3661
timestamp 1714281807
transform 1 0 2848 0 1 370
box -8 -3 16 105
use FILL  FILL_3662
timestamp 1714281807
transform 1 0 2840 0 1 370
box -8 -3 16 105
use FILL  FILL_3663
timestamp 1714281807
transform 1 0 2792 0 1 370
box -8 -3 16 105
use FILL  FILL_3664
timestamp 1714281807
transform 1 0 2784 0 1 370
box -8 -3 16 105
use FILL  FILL_3665
timestamp 1714281807
transform 1 0 2776 0 1 370
box -8 -3 16 105
use FILL  FILL_3666
timestamp 1714281807
transform 1 0 2768 0 1 370
box -8 -3 16 105
use FILL  FILL_3667
timestamp 1714281807
transform 1 0 2760 0 1 370
box -8 -3 16 105
use FILL  FILL_3668
timestamp 1714281807
transform 1 0 2712 0 1 370
box -8 -3 16 105
use FILL  FILL_3669
timestamp 1714281807
transform 1 0 2704 0 1 370
box -8 -3 16 105
use FILL  FILL_3670
timestamp 1714281807
transform 1 0 2696 0 1 370
box -8 -3 16 105
use FILL  FILL_3671
timestamp 1714281807
transform 1 0 2688 0 1 370
box -8 -3 16 105
use FILL  FILL_3672
timestamp 1714281807
transform 1 0 2680 0 1 370
box -8 -3 16 105
use FILL  FILL_3673
timestamp 1714281807
transform 1 0 2584 0 1 370
box -8 -3 16 105
use FILL  FILL_3674
timestamp 1714281807
transform 1 0 2576 0 1 370
box -8 -3 16 105
use FILL  FILL_3675
timestamp 1714281807
transform 1 0 2568 0 1 370
box -8 -3 16 105
use FILL  FILL_3676
timestamp 1714281807
transform 1 0 2520 0 1 370
box -8 -3 16 105
use FILL  FILL_3677
timestamp 1714281807
transform 1 0 2512 0 1 370
box -8 -3 16 105
use FILL  FILL_3678
timestamp 1714281807
transform 1 0 2504 0 1 370
box -8 -3 16 105
use FILL  FILL_3679
timestamp 1714281807
transform 1 0 2496 0 1 370
box -8 -3 16 105
use FILL  FILL_3680
timestamp 1714281807
transform 1 0 2448 0 1 370
box -8 -3 16 105
use FILL  FILL_3681
timestamp 1714281807
transform 1 0 2440 0 1 370
box -8 -3 16 105
use FILL  FILL_3682
timestamp 1714281807
transform 1 0 2432 0 1 370
box -8 -3 16 105
use FILL  FILL_3683
timestamp 1714281807
transform 1 0 2424 0 1 370
box -8 -3 16 105
use FILL  FILL_3684
timestamp 1714281807
transform 1 0 2416 0 1 370
box -8 -3 16 105
use FILL  FILL_3685
timestamp 1714281807
transform 1 0 2408 0 1 370
box -8 -3 16 105
use FILL  FILL_3686
timestamp 1714281807
transform 1 0 2400 0 1 370
box -8 -3 16 105
use FILL  FILL_3687
timestamp 1714281807
transform 1 0 2336 0 1 370
box -8 -3 16 105
use FILL  FILL_3688
timestamp 1714281807
transform 1 0 2328 0 1 370
box -8 -3 16 105
use FILL  FILL_3689
timestamp 1714281807
transform 1 0 2320 0 1 370
box -8 -3 16 105
use FILL  FILL_3690
timestamp 1714281807
transform 1 0 2312 0 1 370
box -8 -3 16 105
use FILL  FILL_3691
timestamp 1714281807
transform 1 0 2304 0 1 370
box -8 -3 16 105
use FILL  FILL_3692
timestamp 1714281807
transform 1 0 2256 0 1 370
box -8 -3 16 105
use FILL  FILL_3693
timestamp 1714281807
transform 1 0 2248 0 1 370
box -8 -3 16 105
use FILL  FILL_3694
timestamp 1714281807
transform 1 0 2240 0 1 370
box -8 -3 16 105
use FILL  FILL_3695
timestamp 1714281807
transform 1 0 2232 0 1 370
box -8 -3 16 105
use FILL  FILL_3696
timestamp 1714281807
transform 1 0 2128 0 1 370
box -8 -3 16 105
use FILL  FILL_3697
timestamp 1714281807
transform 1 0 2120 0 1 370
box -8 -3 16 105
use FILL  FILL_3698
timestamp 1714281807
transform 1 0 2072 0 1 370
box -8 -3 16 105
use FILL  FILL_3699
timestamp 1714281807
transform 1 0 2064 0 1 370
box -8 -3 16 105
use FILL  FILL_3700
timestamp 1714281807
transform 1 0 2056 0 1 370
box -8 -3 16 105
use FILL  FILL_3701
timestamp 1714281807
transform 1 0 2048 0 1 370
box -8 -3 16 105
use FILL  FILL_3702
timestamp 1714281807
transform 1 0 2040 0 1 370
box -8 -3 16 105
use FILL  FILL_3703
timestamp 1714281807
transform 1 0 2032 0 1 370
box -8 -3 16 105
use FILL  FILL_3704
timestamp 1714281807
transform 1 0 1984 0 1 370
box -8 -3 16 105
use FILL  FILL_3705
timestamp 1714281807
transform 1 0 1976 0 1 370
box -8 -3 16 105
use FILL  FILL_3706
timestamp 1714281807
transform 1 0 1968 0 1 370
box -8 -3 16 105
use FILL  FILL_3707
timestamp 1714281807
transform 1 0 1960 0 1 370
box -8 -3 16 105
use FILL  FILL_3708
timestamp 1714281807
transform 1 0 1920 0 1 370
box -8 -3 16 105
use FILL  FILL_3709
timestamp 1714281807
transform 1 0 1912 0 1 370
box -8 -3 16 105
use FILL  FILL_3710
timestamp 1714281807
transform 1 0 1864 0 1 370
box -8 -3 16 105
use FILL  FILL_3711
timestamp 1714281807
transform 1 0 1856 0 1 370
box -8 -3 16 105
use FILL  FILL_3712
timestamp 1714281807
transform 1 0 1848 0 1 370
box -8 -3 16 105
use FILL  FILL_3713
timestamp 1714281807
transform 1 0 1840 0 1 370
box -8 -3 16 105
use FILL  FILL_3714
timestamp 1714281807
transform 1 0 1832 0 1 370
box -8 -3 16 105
use FILL  FILL_3715
timestamp 1714281807
transform 1 0 1824 0 1 370
box -8 -3 16 105
use FILL  FILL_3716
timestamp 1714281807
transform 1 0 1760 0 1 370
box -8 -3 16 105
use FILL  FILL_3717
timestamp 1714281807
transform 1 0 1752 0 1 370
box -8 -3 16 105
use FILL  FILL_3718
timestamp 1714281807
transform 1 0 1744 0 1 370
box -8 -3 16 105
use FILL  FILL_3719
timestamp 1714281807
transform 1 0 1736 0 1 370
box -8 -3 16 105
use FILL  FILL_3720
timestamp 1714281807
transform 1 0 1728 0 1 370
box -8 -3 16 105
use FILL  FILL_3721
timestamp 1714281807
transform 1 0 1680 0 1 370
box -8 -3 16 105
use FILL  FILL_3722
timestamp 1714281807
transform 1 0 1576 0 1 370
box -8 -3 16 105
use FILL  FILL_3723
timestamp 1714281807
transform 1 0 1568 0 1 370
box -8 -3 16 105
use FILL  FILL_3724
timestamp 1714281807
transform 1 0 1520 0 1 370
box -8 -3 16 105
use FILL  FILL_3725
timestamp 1714281807
transform 1 0 1512 0 1 370
box -8 -3 16 105
use FILL  FILL_3726
timestamp 1714281807
transform 1 0 1504 0 1 370
box -8 -3 16 105
use FILL  FILL_3727
timestamp 1714281807
transform 1 0 1496 0 1 370
box -8 -3 16 105
use FILL  FILL_3728
timestamp 1714281807
transform 1 0 1456 0 1 370
box -8 -3 16 105
use FILL  FILL_3729
timestamp 1714281807
transform 1 0 1448 0 1 370
box -8 -3 16 105
use FILL  FILL_3730
timestamp 1714281807
transform 1 0 1400 0 1 370
box -8 -3 16 105
use FILL  FILL_3731
timestamp 1714281807
transform 1 0 1392 0 1 370
box -8 -3 16 105
use FILL  FILL_3732
timestamp 1714281807
transform 1 0 1384 0 1 370
box -8 -3 16 105
use FILL  FILL_3733
timestamp 1714281807
transform 1 0 1320 0 1 370
box -8 -3 16 105
use FILL  FILL_3734
timestamp 1714281807
transform 1 0 1312 0 1 370
box -8 -3 16 105
use FILL  FILL_3735
timestamp 1714281807
transform 1 0 1304 0 1 370
box -8 -3 16 105
use FILL  FILL_3736
timestamp 1714281807
transform 1 0 1256 0 1 370
box -8 -3 16 105
use FILL  FILL_3737
timestamp 1714281807
transform 1 0 1248 0 1 370
box -8 -3 16 105
use FILL  FILL_3738
timestamp 1714281807
transform 1 0 1240 0 1 370
box -8 -3 16 105
use FILL  FILL_3739
timestamp 1714281807
transform 1 0 1232 0 1 370
box -8 -3 16 105
use FILL  FILL_3740
timestamp 1714281807
transform 1 0 1192 0 1 370
box -8 -3 16 105
use FILL  FILL_3741
timestamp 1714281807
transform 1 0 1184 0 1 370
box -8 -3 16 105
use FILL  FILL_3742
timestamp 1714281807
transform 1 0 1176 0 1 370
box -8 -3 16 105
use FILL  FILL_3743
timestamp 1714281807
transform 1 0 1168 0 1 370
box -8 -3 16 105
use FILL  FILL_3744
timestamp 1714281807
transform 1 0 1120 0 1 370
box -8 -3 16 105
use FILL  FILL_3745
timestamp 1714281807
transform 1 0 1112 0 1 370
box -8 -3 16 105
use FILL  FILL_3746
timestamp 1714281807
transform 1 0 1104 0 1 370
box -8 -3 16 105
use FILL  FILL_3747
timestamp 1714281807
transform 1 0 1096 0 1 370
box -8 -3 16 105
use FILL  FILL_3748
timestamp 1714281807
transform 1 0 1088 0 1 370
box -8 -3 16 105
use FILL  FILL_3749
timestamp 1714281807
transform 1 0 1080 0 1 370
box -8 -3 16 105
use FILL  FILL_3750
timestamp 1714281807
transform 1 0 1040 0 1 370
box -8 -3 16 105
use FILL  FILL_3751
timestamp 1714281807
transform 1 0 1016 0 1 370
box -8 -3 16 105
use FILL  FILL_3752
timestamp 1714281807
transform 1 0 1008 0 1 370
box -8 -3 16 105
use FILL  FILL_3753
timestamp 1714281807
transform 1 0 1000 0 1 370
box -8 -3 16 105
use FILL  FILL_3754
timestamp 1714281807
transform 1 0 896 0 1 370
box -8 -3 16 105
use FILL  FILL_3755
timestamp 1714281807
transform 1 0 888 0 1 370
box -8 -3 16 105
use FILL  FILL_3756
timestamp 1714281807
transform 1 0 784 0 1 370
box -8 -3 16 105
use FILL  FILL_3757
timestamp 1714281807
transform 1 0 680 0 1 370
box -8 -3 16 105
use FILL  FILL_3758
timestamp 1714281807
transform 1 0 672 0 1 370
box -8 -3 16 105
use FILL  FILL_3759
timestamp 1714281807
transform 1 0 664 0 1 370
box -8 -3 16 105
use FILL  FILL_3760
timestamp 1714281807
transform 1 0 632 0 1 370
box -8 -3 16 105
use FILL  FILL_3761
timestamp 1714281807
transform 1 0 624 0 1 370
box -8 -3 16 105
use FILL  FILL_3762
timestamp 1714281807
transform 1 0 560 0 1 370
box -8 -3 16 105
use FILL  FILL_3763
timestamp 1714281807
transform 1 0 536 0 1 370
box -8 -3 16 105
use FILL  FILL_3764
timestamp 1714281807
transform 1 0 528 0 1 370
box -8 -3 16 105
use FILL  FILL_3765
timestamp 1714281807
transform 1 0 520 0 1 370
box -8 -3 16 105
use FILL  FILL_3766
timestamp 1714281807
transform 1 0 512 0 1 370
box -8 -3 16 105
use FILL  FILL_3767
timestamp 1714281807
transform 1 0 504 0 1 370
box -8 -3 16 105
use FILL  FILL_3768
timestamp 1714281807
transform 1 0 464 0 1 370
box -8 -3 16 105
use FILL  FILL_3769
timestamp 1714281807
transform 1 0 456 0 1 370
box -8 -3 16 105
use FILL  FILL_3770
timestamp 1714281807
transform 1 0 448 0 1 370
box -8 -3 16 105
use FILL  FILL_3771
timestamp 1714281807
transform 1 0 440 0 1 370
box -8 -3 16 105
use FILL  FILL_3772
timestamp 1714281807
transform 1 0 432 0 1 370
box -8 -3 16 105
use FILL  FILL_3773
timestamp 1714281807
transform 1 0 424 0 1 370
box -8 -3 16 105
use FILL  FILL_3774
timestamp 1714281807
transform 1 0 384 0 1 370
box -8 -3 16 105
use FILL  FILL_3775
timestamp 1714281807
transform 1 0 376 0 1 370
box -8 -3 16 105
use FILL  FILL_3776
timestamp 1714281807
transform 1 0 368 0 1 370
box -8 -3 16 105
use FILL  FILL_3777
timestamp 1714281807
transform 1 0 344 0 1 370
box -8 -3 16 105
use FILL  FILL_3778
timestamp 1714281807
transform 1 0 336 0 1 370
box -8 -3 16 105
use FILL  FILL_3779
timestamp 1714281807
transform 1 0 328 0 1 370
box -8 -3 16 105
use FILL  FILL_3780
timestamp 1714281807
transform 1 0 320 0 1 370
box -8 -3 16 105
use FILL  FILL_3781
timestamp 1714281807
transform 1 0 216 0 1 370
box -8 -3 16 105
use FILL  FILL_3782
timestamp 1714281807
transform 1 0 208 0 1 370
box -8 -3 16 105
use FILL  FILL_3783
timestamp 1714281807
transform 1 0 200 0 1 370
box -8 -3 16 105
use FILL  FILL_3784
timestamp 1714281807
transform 1 0 192 0 1 370
box -8 -3 16 105
use FILL  FILL_3785
timestamp 1714281807
transform 1 0 184 0 1 370
box -8 -3 16 105
use FILL  FILL_3786
timestamp 1714281807
transform 1 0 176 0 1 370
box -8 -3 16 105
use FILL  FILL_3787
timestamp 1714281807
transform 1 0 168 0 1 370
box -8 -3 16 105
use FILL  FILL_3788
timestamp 1714281807
transform 1 0 160 0 1 370
box -8 -3 16 105
use FILL  FILL_3789
timestamp 1714281807
transform 1 0 152 0 1 370
box -8 -3 16 105
use FILL  FILL_3790
timestamp 1714281807
transform 1 0 144 0 1 370
box -8 -3 16 105
use FILL  FILL_3791
timestamp 1714281807
transform 1 0 136 0 1 370
box -8 -3 16 105
use FILL  FILL_3792
timestamp 1714281807
transform 1 0 128 0 1 370
box -8 -3 16 105
use FILL  FILL_3793
timestamp 1714281807
transform 1 0 120 0 1 370
box -8 -3 16 105
use FILL  FILL_3794
timestamp 1714281807
transform 1 0 112 0 1 370
box -8 -3 16 105
use FILL  FILL_3795
timestamp 1714281807
transform 1 0 104 0 1 370
box -8 -3 16 105
use FILL  FILL_3796
timestamp 1714281807
transform 1 0 96 0 1 370
box -8 -3 16 105
use FILL  FILL_3797
timestamp 1714281807
transform 1 0 88 0 1 370
box -8 -3 16 105
use FILL  FILL_3798
timestamp 1714281807
transform 1 0 80 0 1 370
box -8 -3 16 105
use FILL  FILL_3799
timestamp 1714281807
transform 1 0 72 0 1 370
box -8 -3 16 105
use FILL  FILL_3800
timestamp 1714281807
transform 1 0 3000 0 -1 370
box -8 -3 16 105
use FILL  FILL_3801
timestamp 1714281807
transform 1 0 2896 0 -1 370
box -8 -3 16 105
use FILL  FILL_3802
timestamp 1714281807
transform 1 0 2888 0 -1 370
box -8 -3 16 105
use FILL  FILL_3803
timestamp 1714281807
transform 1 0 2864 0 -1 370
box -8 -3 16 105
use FILL  FILL_3804
timestamp 1714281807
transform 1 0 2856 0 -1 370
box -8 -3 16 105
use FILL  FILL_3805
timestamp 1714281807
transform 1 0 2816 0 -1 370
box -8 -3 16 105
use FILL  FILL_3806
timestamp 1714281807
transform 1 0 2808 0 -1 370
box -8 -3 16 105
use FILL  FILL_3807
timestamp 1714281807
transform 1 0 2800 0 -1 370
box -8 -3 16 105
use FILL  FILL_3808
timestamp 1714281807
transform 1 0 2792 0 -1 370
box -8 -3 16 105
use FILL  FILL_3809
timestamp 1714281807
transform 1 0 2784 0 -1 370
box -8 -3 16 105
use FILL  FILL_3810
timestamp 1714281807
transform 1 0 2776 0 -1 370
box -8 -3 16 105
use FILL  FILL_3811
timestamp 1714281807
transform 1 0 2768 0 -1 370
box -8 -3 16 105
use FILL  FILL_3812
timestamp 1714281807
transform 1 0 2728 0 -1 370
box -8 -3 16 105
use FILL  FILL_3813
timestamp 1714281807
transform 1 0 2720 0 -1 370
box -8 -3 16 105
use FILL  FILL_3814
timestamp 1714281807
transform 1 0 2712 0 -1 370
box -8 -3 16 105
use FILL  FILL_3815
timestamp 1714281807
transform 1 0 2704 0 -1 370
box -8 -3 16 105
use FILL  FILL_3816
timestamp 1714281807
transform 1 0 2696 0 -1 370
box -8 -3 16 105
use FILL  FILL_3817
timestamp 1714281807
transform 1 0 2632 0 -1 370
box -8 -3 16 105
use FILL  FILL_3818
timestamp 1714281807
transform 1 0 2624 0 -1 370
box -8 -3 16 105
use FILL  FILL_3819
timestamp 1714281807
transform 1 0 2616 0 -1 370
box -8 -3 16 105
use FILL  FILL_3820
timestamp 1714281807
transform 1 0 2608 0 -1 370
box -8 -3 16 105
use FILL  FILL_3821
timestamp 1714281807
transform 1 0 2600 0 -1 370
box -8 -3 16 105
use FILL  FILL_3822
timestamp 1714281807
transform 1 0 2560 0 -1 370
box -8 -3 16 105
use FILL  FILL_3823
timestamp 1714281807
transform 1 0 2552 0 -1 370
box -8 -3 16 105
use FILL  FILL_3824
timestamp 1714281807
transform 1 0 2544 0 -1 370
box -8 -3 16 105
use FILL  FILL_3825
timestamp 1714281807
transform 1 0 2536 0 -1 370
box -8 -3 16 105
use FILL  FILL_3826
timestamp 1714281807
transform 1 0 2528 0 -1 370
box -8 -3 16 105
use FILL  FILL_3827
timestamp 1714281807
transform 1 0 2520 0 -1 370
box -8 -3 16 105
use FILL  FILL_3828
timestamp 1714281807
transform 1 0 2480 0 -1 370
box -8 -3 16 105
use FILL  FILL_3829
timestamp 1714281807
transform 1 0 2472 0 -1 370
box -8 -3 16 105
use FILL  FILL_3830
timestamp 1714281807
transform 1 0 2464 0 -1 370
box -8 -3 16 105
use FILL  FILL_3831
timestamp 1714281807
transform 1 0 2400 0 -1 370
box -8 -3 16 105
use FILL  FILL_3832
timestamp 1714281807
transform 1 0 2360 0 -1 370
box -8 -3 16 105
use FILL  FILL_3833
timestamp 1714281807
transform 1 0 2352 0 -1 370
box -8 -3 16 105
use FILL  FILL_3834
timestamp 1714281807
transform 1 0 2344 0 -1 370
box -8 -3 16 105
use FILL  FILL_3835
timestamp 1714281807
transform 1 0 2336 0 -1 370
box -8 -3 16 105
use FILL  FILL_3836
timestamp 1714281807
transform 1 0 2328 0 -1 370
box -8 -3 16 105
use FILL  FILL_3837
timestamp 1714281807
transform 1 0 2320 0 -1 370
box -8 -3 16 105
use FILL  FILL_3838
timestamp 1714281807
transform 1 0 2280 0 -1 370
box -8 -3 16 105
use FILL  FILL_3839
timestamp 1714281807
transform 1 0 2272 0 -1 370
box -8 -3 16 105
use FILL  FILL_3840
timestamp 1714281807
transform 1 0 2208 0 -1 370
box -8 -3 16 105
use FILL  FILL_3841
timestamp 1714281807
transform 1 0 2144 0 -1 370
box -8 -3 16 105
use FILL  FILL_3842
timestamp 1714281807
transform 1 0 2136 0 -1 370
box -8 -3 16 105
use FILL  FILL_3843
timestamp 1714281807
transform 1 0 2128 0 -1 370
box -8 -3 16 105
use FILL  FILL_3844
timestamp 1714281807
transform 1 0 2088 0 -1 370
box -8 -3 16 105
use FILL  FILL_3845
timestamp 1714281807
transform 1 0 2080 0 -1 370
box -8 -3 16 105
use FILL  FILL_3846
timestamp 1714281807
transform 1 0 2072 0 -1 370
box -8 -3 16 105
use FILL  FILL_3847
timestamp 1714281807
transform 1 0 2032 0 -1 370
box -8 -3 16 105
use FILL  FILL_3848
timestamp 1714281807
transform 1 0 2024 0 -1 370
box -8 -3 16 105
use FILL  FILL_3849
timestamp 1714281807
transform 1 0 1960 0 -1 370
box -8 -3 16 105
use FILL  FILL_3850
timestamp 1714281807
transform 1 0 1952 0 -1 370
box -8 -3 16 105
use FILL  FILL_3851
timestamp 1714281807
transform 1 0 1912 0 -1 370
box -8 -3 16 105
use FILL  FILL_3852
timestamp 1714281807
transform 1 0 1904 0 -1 370
box -8 -3 16 105
use FILL  FILL_3853
timestamp 1714281807
transform 1 0 1896 0 -1 370
box -8 -3 16 105
use FILL  FILL_3854
timestamp 1714281807
transform 1 0 1888 0 -1 370
box -8 -3 16 105
use FILL  FILL_3855
timestamp 1714281807
transform 1 0 1848 0 -1 370
box -8 -3 16 105
use FILL  FILL_3856
timestamp 1714281807
transform 1 0 1840 0 -1 370
box -8 -3 16 105
use FILL  FILL_3857
timestamp 1714281807
transform 1 0 1720 0 -1 370
box -8 -3 16 105
use FILL  FILL_3858
timestamp 1714281807
transform 1 0 1712 0 -1 370
box -8 -3 16 105
use FILL  FILL_3859
timestamp 1714281807
transform 1 0 1672 0 -1 370
box -8 -3 16 105
use FILL  FILL_3860
timestamp 1714281807
transform 1 0 1664 0 -1 370
box -8 -3 16 105
use FILL  FILL_3861
timestamp 1714281807
transform 1 0 1656 0 -1 370
box -8 -3 16 105
use FILL  FILL_3862
timestamp 1714281807
transform 1 0 1648 0 -1 370
box -8 -3 16 105
use FILL  FILL_3863
timestamp 1714281807
transform 1 0 1608 0 -1 370
box -8 -3 16 105
use FILL  FILL_3864
timestamp 1714281807
transform 1 0 1600 0 -1 370
box -8 -3 16 105
use FILL  FILL_3865
timestamp 1714281807
transform 1 0 1592 0 -1 370
box -8 -3 16 105
use FILL  FILL_3866
timestamp 1714281807
transform 1 0 1528 0 -1 370
box -8 -3 16 105
use FILL  FILL_3867
timestamp 1714281807
transform 1 0 1488 0 -1 370
box -8 -3 16 105
use FILL  FILL_3868
timestamp 1714281807
transform 1 0 1480 0 -1 370
box -8 -3 16 105
use FILL  FILL_3869
timestamp 1714281807
transform 1 0 1472 0 -1 370
box -8 -3 16 105
use FILL  FILL_3870
timestamp 1714281807
transform 1 0 1464 0 -1 370
box -8 -3 16 105
use FILL  FILL_3871
timestamp 1714281807
transform 1 0 1456 0 -1 370
box -8 -3 16 105
use FILL  FILL_3872
timestamp 1714281807
transform 1 0 1448 0 -1 370
box -8 -3 16 105
use FILL  FILL_3873
timestamp 1714281807
transform 1 0 1440 0 -1 370
box -8 -3 16 105
use FILL  FILL_3874
timestamp 1714281807
transform 1 0 1400 0 -1 370
box -8 -3 16 105
use FILL  FILL_3875
timestamp 1714281807
transform 1 0 1392 0 -1 370
box -8 -3 16 105
use FILL  FILL_3876
timestamp 1714281807
transform 1 0 1384 0 -1 370
box -8 -3 16 105
use FILL  FILL_3877
timestamp 1714281807
transform 1 0 1376 0 -1 370
box -8 -3 16 105
use FILL  FILL_3878
timestamp 1714281807
transform 1 0 1312 0 -1 370
box -8 -3 16 105
use FILL  FILL_3879
timestamp 1714281807
transform 1 0 1304 0 -1 370
box -8 -3 16 105
use FILL  FILL_3880
timestamp 1714281807
transform 1 0 1296 0 -1 370
box -8 -3 16 105
use FILL  FILL_3881
timestamp 1714281807
transform 1 0 1256 0 -1 370
box -8 -3 16 105
use FILL  FILL_3882
timestamp 1714281807
transform 1 0 1248 0 -1 370
box -8 -3 16 105
use FILL  FILL_3883
timestamp 1714281807
transform 1 0 1240 0 -1 370
box -8 -3 16 105
use FILL  FILL_3884
timestamp 1714281807
transform 1 0 1232 0 -1 370
box -8 -3 16 105
use FILL  FILL_3885
timestamp 1714281807
transform 1 0 1224 0 -1 370
box -8 -3 16 105
use FILL  FILL_3886
timestamp 1714281807
transform 1 0 1216 0 -1 370
box -8 -3 16 105
use FILL  FILL_3887
timestamp 1714281807
transform 1 0 1168 0 -1 370
box -8 -3 16 105
use FILL  FILL_3888
timestamp 1714281807
transform 1 0 1160 0 -1 370
box -8 -3 16 105
use FILL  FILL_3889
timestamp 1714281807
transform 1 0 1152 0 -1 370
box -8 -3 16 105
use FILL  FILL_3890
timestamp 1714281807
transform 1 0 1144 0 -1 370
box -8 -3 16 105
use FILL  FILL_3891
timestamp 1714281807
transform 1 0 1136 0 -1 370
box -8 -3 16 105
use FILL  FILL_3892
timestamp 1714281807
transform 1 0 1128 0 -1 370
box -8 -3 16 105
use FILL  FILL_3893
timestamp 1714281807
transform 1 0 1088 0 -1 370
box -8 -3 16 105
use FILL  FILL_3894
timestamp 1714281807
transform 1 0 1080 0 -1 370
box -8 -3 16 105
use FILL  FILL_3895
timestamp 1714281807
transform 1 0 1072 0 -1 370
box -8 -3 16 105
use FILL  FILL_3896
timestamp 1714281807
transform 1 0 1064 0 -1 370
box -8 -3 16 105
use FILL  FILL_3897
timestamp 1714281807
transform 1 0 1056 0 -1 370
box -8 -3 16 105
use FILL  FILL_3898
timestamp 1714281807
transform 1 0 1024 0 -1 370
box -8 -3 16 105
use FILL  FILL_3899
timestamp 1714281807
transform 1 0 1016 0 -1 370
box -8 -3 16 105
use FILL  FILL_3900
timestamp 1714281807
transform 1 0 1008 0 -1 370
box -8 -3 16 105
use FILL  FILL_3901
timestamp 1714281807
transform 1 0 904 0 -1 370
box -8 -3 16 105
use FILL  FILL_3902
timestamp 1714281807
transform 1 0 896 0 -1 370
box -8 -3 16 105
use FILL  FILL_3903
timestamp 1714281807
transform 1 0 888 0 -1 370
box -8 -3 16 105
use FILL  FILL_3904
timestamp 1714281807
transform 1 0 864 0 -1 370
box -8 -3 16 105
use FILL  FILL_3905
timestamp 1714281807
transform 1 0 856 0 -1 370
box -8 -3 16 105
use FILL  FILL_3906
timestamp 1714281807
transform 1 0 848 0 -1 370
box -8 -3 16 105
use FILL  FILL_3907
timestamp 1714281807
transform 1 0 816 0 -1 370
box -8 -3 16 105
use FILL  FILL_3908
timestamp 1714281807
transform 1 0 808 0 -1 370
box -8 -3 16 105
use FILL  FILL_3909
timestamp 1714281807
transform 1 0 800 0 -1 370
box -8 -3 16 105
use FILL  FILL_3910
timestamp 1714281807
transform 1 0 792 0 -1 370
box -8 -3 16 105
use FILL  FILL_3911
timestamp 1714281807
transform 1 0 784 0 -1 370
box -8 -3 16 105
use FILL  FILL_3912
timestamp 1714281807
transform 1 0 744 0 -1 370
box -8 -3 16 105
use FILL  FILL_3913
timestamp 1714281807
transform 1 0 736 0 -1 370
box -8 -3 16 105
use FILL  FILL_3914
timestamp 1714281807
transform 1 0 728 0 -1 370
box -8 -3 16 105
use FILL  FILL_3915
timestamp 1714281807
transform 1 0 720 0 -1 370
box -8 -3 16 105
use FILL  FILL_3916
timestamp 1714281807
transform 1 0 712 0 -1 370
box -8 -3 16 105
use FILL  FILL_3917
timestamp 1714281807
transform 1 0 672 0 -1 370
box -8 -3 16 105
use FILL  FILL_3918
timestamp 1714281807
transform 1 0 664 0 -1 370
box -8 -3 16 105
use FILL  FILL_3919
timestamp 1714281807
transform 1 0 656 0 -1 370
box -8 -3 16 105
use FILL  FILL_3920
timestamp 1714281807
transform 1 0 616 0 -1 370
box -8 -3 16 105
use FILL  FILL_3921
timestamp 1714281807
transform 1 0 608 0 -1 370
box -8 -3 16 105
use FILL  FILL_3922
timestamp 1714281807
transform 1 0 600 0 -1 370
box -8 -3 16 105
use FILL  FILL_3923
timestamp 1714281807
transform 1 0 592 0 -1 370
box -8 -3 16 105
use FILL  FILL_3924
timestamp 1714281807
transform 1 0 584 0 -1 370
box -8 -3 16 105
use FILL  FILL_3925
timestamp 1714281807
transform 1 0 544 0 -1 370
box -8 -3 16 105
use FILL  FILL_3926
timestamp 1714281807
transform 1 0 536 0 -1 370
box -8 -3 16 105
use FILL  FILL_3927
timestamp 1714281807
transform 1 0 528 0 -1 370
box -8 -3 16 105
use FILL  FILL_3928
timestamp 1714281807
transform 1 0 520 0 -1 370
box -8 -3 16 105
use FILL  FILL_3929
timestamp 1714281807
transform 1 0 472 0 -1 370
box -8 -3 16 105
use FILL  FILL_3930
timestamp 1714281807
transform 1 0 464 0 -1 370
box -8 -3 16 105
use FILL  FILL_3931
timestamp 1714281807
transform 1 0 456 0 -1 370
box -8 -3 16 105
use FILL  FILL_3932
timestamp 1714281807
transform 1 0 448 0 -1 370
box -8 -3 16 105
use FILL  FILL_3933
timestamp 1714281807
transform 1 0 440 0 -1 370
box -8 -3 16 105
use FILL  FILL_3934
timestamp 1714281807
transform 1 0 432 0 -1 370
box -8 -3 16 105
use FILL  FILL_3935
timestamp 1714281807
transform 1 0 392 0 -1 370
box -8 -3 16 105
use FILL  FILL_3936
timestamp 1714281807
transform 1 0 368 0 -1 370
box -8 -3 16 105
use FILL  FILL_3937
timestamp 1714281807
transform 1 0 360 0 -1 370
box -8 -3 16 105
use FILL  FILL_3938
timestamp 1714281807
transform 1 0 352 0 -1 370
box -8 -3 16 105
use FILL  FILL_3939
timestamp 1714281807
transform 1 0 344 0 -1 370
box -8 -3 16 105
use FILL  FILL_3940
timestamp 1714281807
transform 1 0 336 0 -1 370
box -8 -3 16 105
use FILL  FILL_3941
timestamp 1714281807
transform 1 0 328 0 -1 370
box -8 -3 16 105
use FILL  FILL_3942
timestamp 1714281807
transform 1 0 280 0 -1 370
box -8 -3 16 105
use FILL  FILL_3943
timestamp 1714281807
transform 1 0 272 0 -1 370
box -8 -3 16 105
use FILL  FILL_3944
timestamp 1714281807
transform 1 0 264 0 -1 370
box -8 -3 16 105
use FILL  FILL_3945
timestamp 1714281807
transform 1 0 256 0 -1 370
box -8 -3 16 105
use FILL  FILL_3946
timestamp 1714281807
transform 1 0 248 0 -1 370
box -8 -3 16 105
use FILL  FILL_3947
timestamp 1714281807
transform 1 0 240 0 -1 370
box -8 -3 16 105
use FILL  FILL_3948
timestamp 1714281807
transform 1 0 208 0 -1 370
box -8 -3 16 105
use FILL  FILL_3949
timestamp 1714281807
transform 1 0 200 0 -1 370
box -8 -3 16 105
use FILL  FILL_3950
timestamp 1714281807
transform 1 0 192 0 -1 370
box -8 -3 16 105
use FILL  FILL_3951
timestamp 1714281807
transform 1 0 184 0 -1 370
box -8 -3 16 105
use FILL  FILL_3952
timestamp 1714281807
transform 1 0 176 0 -1 370
box -8 -3 16 105
use FILL  FILL_3953
timestamp 1714281807
transform 1 0 168 0 -1 370
box -8 -3 16 105
use FILL  FILL_3954
timestamp 1714281807
transform 1 0 160 0 -1 370
box -8 -3 16 105
use FILL  FILL_3955
timestamp 1714281807
transform 1 0 152 0 -1 370
box -8 -3 16 105
use FILL  FILL_3956
timestamp 1714281807
transform 1 0 144 0 -1 370
box -8 -3 16 105
use FILL  FILL_3957
timestamp 1714281807
transform 1 0 136 0 -1 370
box -8 -3 16 105
use FILL  FILL_3958
timestamp 1714281807
transform 1 0 128 0 -1 370
box -8 -3 16 105
use FILL  FILL_3959
timestamp 1714281807
transform 1 0 120 0 -1 370
box -8 -3 16 105
use FILL  FILL_3960
timestamp 1714281807
transform 1 0 112 0 -1 370
box -8 -3 16 105
use FILL  FILL_3961
timestamp 1714281807
transform 1 0 104 0 -1 370
box -8 -3 16 105
use FILL  FILL_3962
timestamp 1714281807
transform 1 0 96 0 -1 370
box -8 -3 16 105
use FILL  FILL_3963
timestamp 1714281807
transform 1 0 88 0 -1 370
box -8 -3 16 105
use FILL  FILL_3964
timestamp 1714281807
transform 1 0 80 0 -1 370
box -8 -3 16 105
use FILL  FILL_3965
timestamp 1714281807
transform 1 0 72 0 -1 370
box -8 -3 16 105
use FILL  FILL_3966
timestamp 1714281807
transform 1 0 3000 0 1 170
box -8 -3 16 105
use FILL  FILL_3967
timestamp 1714281807
transform 1 0 2896 0 1 170
box -8 -3 16 105
use FILL  FILL_3968
timestamp 1714281807
transform 1 0 2888 0 1 170
box -8 -3 16 105
use FILL  FILL_3969
timestamp 1714281807
transform 1 0 2880 0 1 170
box -8 -3 16 105
use FILL  FILL_3970
timestamp 1714281807
transform 1 0 2872 0 1 170
box -8 -3 16 105
use FILL  FILL_3971
timestamp 1714281807
transform 1 0 2840 0 1 170
box -8 -3 16 105
use FILL  FILL_3972
timestamp 1714281807
transform 1 0 2832 0 1 170
box -8 -3 16 105
use FILL  FILL_3973
timestamp 1714281807
transform 1 0 2824 0 1 170
box -8 -3 16 105
use FILL  FILL_3974
timestamp 1714281807
transform 1 0 2816 0 1 170
box -8 -3 16 105
use FILL  FILL_3975
timestamp 1714281807
transform 1 0 2808 0 1 170
box -8 -3 16 105
use FILL  FILL_3976
timestamp 1714281807
transform 1 0 2704 0 1 170
box -8 -3 16 105
use FILL  FILL_3977
timestamp 1714281807
transform 1 0 2680 0 1 170
box -8 -3 16 105
use FILL  FILL_3978
timestamp 1714281807
transform 1 0 2672 0 1 170
box -8 -3 16 105
use FILL  FILL_3979
timestamp 1714281807
transform 1 0 2664 0 1 170
box -8 -3 16 105
use FILL  FILL_3980
timestamp 1714281807
transform 1 0 2656 0 1 170
box -8 -3 16 105
use FILL  FILL_3981
timestamp 1714281807
transform 1 0 2648 0 1 170
box -8 -3 16 105
use FILL  FILL_3982
timestamp 1714281807
transform 1 0 2640 0 1 170
box -8 -3 16 105
use FILL  FILL_3983
timestamp 1714281807
transform 1 0 2424 0 1 170
box -8 -3 16 105
use FILL  FILL_3984
timestamp 1714281807
transform 1 0 2400 0 1 170
box -8 -3 16 105
use FILL  FILL_3985
timestamp 1714281807
transform 1 0 2392 0 1 170
box -8 -3 16 105
use FILL  FILL_3986
timestamp 1714281807
transform 1 0 2384 0 1 170
box -8 -3 16 105
use FILL  FILL_3987
timestamp 1714281807
transform 1 0 2376 0 1 170
box -8 -3 16 105
use FILL  FILL_3988
timestamp 1714281807
transform 1 0 2368 0 1 170
box -8 -3 16 105
use FILL  FILL_3989
timestamp 1714281807
transform 1 0 2360 0 1 170
box -8 -3 16 105
use FILL  FILL_3990
timestamp 1714281807
transform 1 0 2352 0 1 170
box -8 -3 16 105
use FILL  FILL_3991
timestamp 1714281807
transform 1 0 2232 0 1 170
box -8 -3 16 105
use FILL  FILL_3992
timestamp 1714281807
transform 1 0 2224 0 1 170
box -8 -3 16 105
use FILL  FILL_3993
timestamp 1714281807
transform 1 0 2216 0 1 170
box -8 -3 16 105
use FILL  FILL_3994
timestamp 1714281807
transform 1 0 2112 0 1 170
box -8 -3 16 105
use FILL  FILL_3995
timestamp 1714281807
transform 1 0 2104 0 1 170
box -8 -3 16 105
use FILL  FILL_3996
timestamp 1714281807
transform 1 0 2080 0 1 170
box -8 -3 16 105
use FILL  FILL_3997
timestamp 1714281807
transform 1 0 2056 0 1 170
box -8 -3 16 105
use FILL  FILL_3998
timestamp 1714281807
transform 1 0 2048 0 1 170
box -8 -3 16 105
use FILL  FILL_3999
timestamp 1714281807
transform 1 0 1944 0 1 170
box -8 -3 16 105
use FILL  FILL_4000
timestamp 1714281807
transform 1 0 1936 0 1 170
box -8 -3 16 105
use FILL  FILL_4001
timestamp 1714281807
transform 1 0 1832 0 1 170
box -8 -3 16 105
use FILL  FILL_4002
timestamp 1714281807
transform 1 0 1824 0 1 170
box -8 -3 16 105
use FILL  FILL_4003
timestamp 1714281807
transform 1 0 1800 0 1 170
box -8 -3 16 105
use FILL  FILL_4004
timestamp 1714281807
transform 1 0 1792 0 1 170
box -8 -3 16 105
use FILL  FILL_4005
timestamp 1714281807
transform 1 0 1784 0 1 170
box -8 -3 16 105
use FILL  FILL_4006
timestamp 1714281807
transform 1 0 1776 0 1 170
box -8 -3 16 105
use FILL  FILL_4007
timestamp 1714281807
transform 1 0 1768 0 1 170
box -8 -3 16 105
use FILL  FILL_4008
timestamp 1714281807
transform 1 0 1744 0 1 170
box -8 -3 16 105
use FILL  FILL_4009
timestamp 1714281807
transform 1 0 1736 0 1 170
box -8 -3 16 105
use FILL  FILL_4010
timestamp 1714281807
transform 1 0 1632 0 1 170
box -8 -3 16 105
use FILL  FILL_4011
timestamp 1714281807
transform 1 0 1624 0 1 170
box -8 -3 16 105
use FILL  FILL_4012
timestamp 1714281807
transform 1 0 1616 0 1 170
box -8 -3 16 105
use FILL  FILL_4013
timestamp 1714281807
transform 1 0 1496 0 1 170
box -8 -3 16 105
use FILL  FILL_4014
timestamp 1714281807
transform 1 0 1488 0 1 170
box -8 -3 16 105
use FILL  FILL_4015
timestamp 1714281807
transform 1 0 1480 0 1 170
box -8 -3 16 105
use FILL  FILL_4016
timestamp 1714281807
transform 1 0 1472 0 1 170
box -8 -3 16 105
use FILL  FILL_4017
timestamp 1714281807
transform 1 0 1352 0 1 170
box -8 -3 16 105
use FILL  FILL_4018
timestamp 1714281807
transform 1 0 1344 0 1 170
box -8 -3 16 105
use FILL  FILL_4019
timestamp 1714281807
transform 1 0 1336 0 1 170
box -8 -3 16 105
use FILL  FILL_4020
timestamp 1714281807
transform 1 0 1232 0 1 170
box -8 -3 16 105
use FILL  FILL_4021
timestamp 1714281807
transform 1 0 1224 0 1 170
box -8 -3 16 105
use FILL  FILL_4022
timestamp 1714281807
transform 1 0 1200 0 1 170
box -8 -3 16 105
use FILL  FILL_4023
timestamp 1714281807
transform 1 0 1192 0 1 170
box -8 -3 16 105
use FILL  FILL_4024
timestamp 1714281807
transform 1 0 1184 0 1 170
box -8 -3 16 105
use FILL  FILL_4025
timestamp 1714281807
transform 1 0 1160 0 1 170
box -8 -3 16 105
use FILL  FILL_4026
timestamp 1714281807
transform 1 0 1152 0 1 170
box -8 -3 16 105
use FILL  FILL_4027
timestamp 1714281807
transform 1 0 1048 0 1 170
box -8 -3 16 105
use FILL  FILL_4028
timestamp 1714281807
transform 1 0 1040 0 1 170
box -8 -3 16 105
use FILL  FILL_4029
timestamp 1714281807
transform 1 0 1032 0 1 170
box -8 -3 16 105
use FILL  FILL_4030
timestamp 1714281807
transform 1 0 1024 0 1 170
box -8 -3 16 105
use FILL  FILL_4031
timestamp 1714281807
transform 1 0 1016 0 1 170
box -8 -3 16 105
use FILL  FILL_4032
timestamp 1714281807
transform 1 0 984 0 1 170
box -8 -3 16 105
use FILL  FILL_4033
timestamp 1714281807
transform 1 0 976 0 1 170
box -8 -3 16 105
use FILL  FILL_4034
timestamp 1714281807
transform 1 0 968 0 1 170
box -8 -3 16 105
use FILL  FILL_4035
timestamp 1714281807
transform 1 0 960 0 1 170
box -8 -3 16 105
use FILL  FILL_4036
timestamp 1714281807
transform 1 0 952 0 1 170
box -8 -3 16 105
use FILL  FILL_4037
timestamp 1714281807
transform 1 0 944 0 1 170
box -8 -3 16 105
use FILL  FILL_4038
timestamp 1714281807
transform 1 0 936 0 1 170
box -8 -3 16 105
use FILL  FILL_4039
timestamp 1714281807
transform 1 0 928 0 1 170
box -8 -3 16 105
use FILL  FILL_4040
timestamp 1714281807
transform 1 0 920 0 1 170
box -8 -3 16 105
use FILL  FILL_4041
timestamp 1714281807
transform 1 0 912 0 1 170
box -8 -3 16 105
use FILL  FILL_4042
timestamp 1714281807
transform 1 0 904 0 1 170
box -8 -3 16 105
use FILL  FILL_4043
timestamp 1714281807
transform 1 0 896 0 1 170
box -8 -3 16 105
use FILL  FILL_4044
timestamp 1714281807
transform 1 0 888 0 1 170
box -8 -3 16 105
use FILL  FILL_4045
timestamp 1714281807
transform 1 0 880 0 1 170
box -8 -3 16 105
use FILL  FILL_4046
timestamp 1714281807
transform 1 0 872 0 1 170
box -8 -3 16 105
use FILL  FILL_4047
timestamp 1714281807
transform 1 0 864 0 1 170
box -8 -3 16 105
use FILL  FILL_4048
timestamp 1714281807
transform 1 0 856 0 1 170
box -8 -3 16 105
use FILL  FILL_4049
timestamp 1714281807
transform 1 0 848 0 1 170
box -8 -3 16 105
use FILL  FILL_4050
timestamp 1714281807
transform 1 0 840 0 1 170
box -8 -3 16 105
use FILL  FILL_4051
timestamp 1714281807
transform 1 0 832 0 1 170
box -8 -3 16 105
use FILL  FILL_4052
timestamp 1714281807
transform 1 0 824 0 1 170
box -8 -3 16 105
use FILL  FILL_4053
timestamp 1714281807
transform 1 0 816 0 1 170
box -8 -3 16 105
use FILL  FILL_4054
timestamp 1714281807
transform 1 0 808 0 1 170
box -8 -3 16 105
use FILL  FILL_4055
timestamp 1714281807
transform 1 0 800 0 1 170
box -8 -3 16 105
use FILL  FILL_4056
timestamp 1714281807
transform 1 0 792 0 1 170
box -8 -3 16 105
use FILL  FILL_4057
timestamp 1714281807
transform 1 0 784 0 1 170
box -8 -3 16 105
use FILL  FILL_4058
timestamp 1714281807
transform 1 0 776 0 1 170
box -8 -3 16 105
use FILL  FILL_4059
timestamp 1714281807
transform 1 0 736 0 1 170
box -8 -3 16 105
use FILL  FILL_4060
timestamp 1714281807
transform 1 0 728 0 1 170
box -8 -3 16 105
use FILL  FILL_4061
timestamp 1714281807
transform 1 0 720 0 1 170
box -8 -3 16 105
use FILL  FILL_4062
timestamp 1714281807
transform 1 0 712 0 1 170
box -8 -3 16 105
use FILL  FILL_4063
timestamp 1714281807
transform 1 0 704 0 1 170
box -8 -3 16 105
use FILL  FILL_4064
timestamp 1714281807
transform 1 0 696 0 1 170
box -8 -3 16 105
use FILL  FILL_4065
timestamp 1714281807
transform 1 0 688 0 1 170
box -8 -3 16 105
use FILL  FILL_4066
timestamp 1714281807
transform 1 0 664 0 1 170
box -8 -3 16 105
use FILL  FILL_4067
timestamp 1714281807
transform 1 0 656 0 1 170
box -8 -3 16 105
use FILL  FILL_4068
timestamp 1714281807
transform 1 0 632 0 1 170
box -8 -3 16 105
use FILL  FILL_4069
timestamp 1714281807
transform 1 0 624 0 1 170
box -8 -3 16 105
use FILL  FILL_4070
timestamp 1714281807
transform 1 0 616 0 1 170
box -8 -3 16 105
use FILL  FILL_4071
timestamp 1714281807
transform 1 0 608 0 1 170
box -8 -3 16 105
use FILL  FILL_4072
timestamp 1714281807
transform 1 0 600 0 1 170
box -8 -3 16 105
use FILL  FILL_4073
timestamp 1714281807
transform 1 0 592 0 1 170
box -8 -3 16 105
use FILL  FILL_4074
timestamp 1714281807
transform 1 0 560 0 1 170
box -8 -3 16 105
use FILL  FILL_4075
timestamp 1714281807
transform 1 0 552 0 1 170
box -8 -3 16 105
use FILL  FILL_4076
timestamp 1714281807
transform 1 0 544 0 1 170
box -8 -3 16 105
use FILL  FILL_4077
timestamp 1714281807
transform 1 0 536 0 1 170
box -8 -3 16 105
use FILL  FILL_4078
timestamp 1714281807
transform 1 0 528 0 1 170
box -8 -3 16 105
use FILL  FILL_4079
timestamp 1714281807
transform 1 0 520 0 1 170
box -8 -3 16 105
use FILL  FILL_4080
timestamp 1714281807
transform 1 0 480 0 1 170
box -8 -3 16 105
use FILL  FILL_4081
timestamp 1714281807
transform 1 0 472 0 1 170
box -8 -3 16 105
use FILL  FILL_4082
timestamp 1714281807
transform 1 0 464 0 1 170
box -8 -3 16 105
use FILL  FILL_4083
timestamp 1714281807
transform 1 0 456 0 1 170
box -8 -3 16 105
use FILL  FILL_4084
timestamp 1714281807
transform 1 0 448 0 1 170
box -8 -3 16 105
use FILL  FILL_4085
timestamp 1714281807
transform 1 0 440 0 1 170
box -8 -3 16 105
use FILL  FILL_4086
timestamp 1714281807
transform 1 0 416 0 1 170
box -8 -3 16 105
use FILL  FILL_4087
timestamp 1714281807
transform 1 0 408 0 1 170
box -8 -3 16 105
use FILL  FILL_4088
timestamp 1714281807
transform 1 0 400 0 1 170
box -8 -3 16 105
use FILL  FILL_4089
timestamp 1714281807
transform 1 0 392 0 1 170
box -8 -3 16 105
use FILL  FILL_4090
timestamp 1714281807
transform 1 0 352 0 1 170
box -8 -3 16 105
use FILL  FILL_4091
timestamp 1714281807
transform 1 0 344 0 1 170
box -8 -3 16 105
use FILL  FILL_4092
timestamp 1714281807
transform 1 0 336 0 1 170
box -8 -3 16 105
use FILL  FILL_4093
timestamp 1714281807
transform 1 0 328 0 1 170
box -8 -3 16 105
use FILL  FILL_4094
timestamp 1714281807
transform 1 0 320 0 1 170
box -8 -3 16 105
use FILL  FILL_4095
timestamp 1714281807
transform 1 0 312 0 1 170
box -8 -3 16 105
use FILL  FILL_4096
timestamp 1714281807
transform 1 0 304 0 1 170
box -8 -3 16 105
use FILL  FILL_4097
timestamp 1714281807
transform 1 0 272 0 1 170
box -8 -3 16 105
use FILL  FILL_4098
timestamp 1714281807
transform 1 0 264 0 1 170
box -8 -3 16 105
use FILL  FILL_4099
timestamp 1714281807
transform 1 0 256 0 1 170
box -8 -3 16 105
use FILL  FILL_4100
timestamp 1714281807
transform 1 0 248 0 1 170
box -8 -3 16 105
use FILL  FILL_4101
timestamp 1714281807
transform 1 0 240 0 1 170
box -8 -3 16 105
use FILL  FILL_4102
timestamp 1714281807
transform 1 0 232 0 1 170
box -8 -3 16 105
use FILL  FILL_4103
timestamp 1714281807
transform 1 0 224 0 1 170
box -8 -3 16 105
use FILL  FILL_4104
timestamp 1714281807
transform 1 0 216 0 1 170
box -8 -3 16 105
use FILL  FILL_4105
timestamp 1714281807
transform 1 0 208 0 1 170
box -8 -3 16 105
use FILL  FILL_4106
timestamp 1714281807
transform 1 0 200 0 1 170
box -8 -3 16 105
use FILL  FILL_4107
timestamp 1714281807
transform 1 0 192 0 1 170
box -8 -3 16 105
use FILL  FILL_4108
timestamp 1714281807
transform 1 0 184 0 1 170
box -8 -3 16 105
use FILL  FILL_4109
timestamp 1714281807
transform 1 0 176 0 1 170
box -8 -3 16 105
use FILL  FILL_4110
timestamp 1714281807
transform 1 0 168 0 1 170
box -8 -3 16 105
use FILL  FILL_4111
timestamp 1714281807
transform 1 0 160 0 1 170
box -8 -3 16 105
use FILL  FILL_4112
timestamp 1714281807
transform 1 0 152 0 1 170
box -8 -3 16 105
use FILL  FILL_4113
timestamp 1714281807
transform 1 0 144 0 1 170
box -8 -3 16 105
use FILL  FILL_4114
timestamp 1714281807
transform 1 0 136 0 1 170
box -8 -3 16 105
use FILL  FILL_4115
timestamp 1714281807
transform 1 0 128 0 1 170
box -8 -3 16 105
use FILL  FILL_4116
timestamp 1714281807
transform 1 0 120 0 1 170
box -8 -3 16 105
use FILL  FILL_4117
timestamp 1714281807
transform 1 0 112 0 1 170
box -8 -3 16 105
use FILL  FILL_4118
timestamp 1714281807
transform 1 0 104 0 1 170
box -8 -3 16 105
use FILL  FILL_4119
timestamp 1714281807
transform 1 0 96 0 1 170
box -8 -3 16 105
use FILL  FILL_4120
timestamp 1714281807
transform 1 0 88 0 1 170
box -8 -3 16 105
use FILL  FILL_4121
timestamp 1714281807
transform 1 0 80 0 1 170
box -8 -3 16 105
use FILL  FILL_4122
timestamp 1714281807
transform 1 0 72 0 1 170
box -8 -3 16 105
use FILL  FILL_4123
timestamp 1714281807
transform 1 0 3000 0 -1 170
box -8 -3 16 105
use FILL  FILL_4124
timestamp 1714281807
transform 1 0 2896 0 -1 170
box -8 -3 16 105
use FILL  FILL_4125
timestamp 1714281807
transform 1 0 2888 0 -1 170
box -8 -3 16 105
use FILL  FILL_4126
timestamp 1714281807
transform 1 0 2856 0 -1 170
box -8 -3 16 105
use FILL  FILL_4127
timestamp 1714281807
transform 1 0 2848 0 -1 170
box -8 -3 16 105
use FILL  FILL_4128
timestamp 1714281807
transform 1 0 2720 0 -1 170
box -8 -3 16 105
use FILL  FILL_4129
timestamp 1714281807
transform 1 0 2712 0 -1 170
box -8 -3 16 105
use FILL  FILL_4130
timestamp 1714281807
transform 1 0 2608 0 -1 170
box -8 -3 16 105
use FILL  FILL_4131
timestamp 1714281807
transform 1 0 2576 0 -1 170
box -8 -3 16 105
use FILL  FILL_4132
timestamp 1714281807
transform 1 0 2568 0 -1 170
box -8 -3 16 105
use FILL  FILL_4133
timestamp 1714281807
transform 1 0 2464 0 -1 170
box -8 -3 16 105
use FILL  FILL_4134
timestamp 1714281807
transform 1 0 2456 0 -1 170
box -8 -3 16 105
use FILL  FILL_4135
timestamp 1714281807
transform 1 0 2448 0 -1 170
box -8 -3 16 105
use FILL  FILL_4136
timestamp 1714281807
transform 1 0 2416 0 -1 170
box -8 -3 16 105
use FILL  FILL_4137
timestamp 1714281807
transform 1 0 2408 0 -1 170
box -8 -3 16 105
use FILL  FILL_4138
timestamp 1714281807
transform 1 0 2400 0 -1 170
box -8 -3 16 105
use FILL  FILL_4139
timestamp 1714281807
transform 1 0 2392 0 -1 170
box -8 -3 16 105
use FILL  FILL_4140
timestamp 1714281807
transform 1 0 2288 0 -1 170
box -8 -3 16 105
use FILL  FILL_4141
timestamp 1714281807
transform 1 0 2280 0 -1 170
box -8 -3 16 105
use FILL  FILL_4142
timestamp 1714281807
transform 1 0 2272 0 -1 170
box -8 -3 16 105
use FILL  FILL_4143
timestamp 1714281807
transform 1 0 2240 0 -1 170
box -8 -3 16 105
use FILL  FILL_4144
timestamp 1714281807
transform 1 0 2232 0 -1 170
box -8 -3 16 105
use FILL  FILL_4145
timestamp 1714281807
transform 1 0 2224 0 -1 170
box -8 -3 16 105
use FILL  FILL_4146
timestamp 1714281807
transform 1 0 2216 0 -1 170
box -8 -3 16 105
use FILL  FILL_4147
timestamp 1714281807
transform 1 0 2112 0 -1 170
box -8 -3 16 105
use FILL  FILL_4148
timestamp 1714281807
transform 1 0 2104 0 -1 170
box -8 -3 16 105
use FILL  FILL_4149
timestamp 1714281807
transform 1 0 2096 0 -1 170
box -8 -3 16 105
use FILL  FILL_4150
timestamp 1714281807
transform 1 0 2088 0 -1 170
box -8 -3 16 105
use FILL  FILL_4151
timestamp 1714281807
transform 1 0 2056 0 -1 170
box -8 -3 16 105
use FILL  FILL_4152
timestamp 1714281807
transform 1 0 2048 0 -1 170
box -8 -3 16 105
use FILL  FILL_4153
timestamp 1714281807
transform 1 0 2040 0 -1 170
box -8 -3 16 105
use FILL  FILL_4154
timestamp 1714281807
transform 1 0 2008 0 -1 170
box -8 -3 16 105
use FILL  FILL_4155
timestamp 1714281807
transform 1 0 2000 0 -1 170
box -8 -3 16 105
use FILL  FILL_4156
timestamp 1714281807
transform 1 0 1992 0 -1 170
box -8 -3 16 105
use FILL  FILL_4157
timestamp 1714281807
transform 1 0 1984 0 -1 170
box -8 -3 16 105
use FILL  FILL_4158
timestamp 1714281807
transform 1 0 1880 0 -1 170
box -8 -3 16 105
use FILL  FILL_4159
timestamp 1714281807
transform 1 0 1872 0 -1 170
box -8 -3 16 105
use FILL  FILL_4160
timestamp 1714281807
transform 1 0 1840 0 -1 170
box -8 -3 16 105
use FILL  FILL_4161
timestamp 1714281807
transform 1 0 1832 0 -1 170
box -8 -3 16 105
use FILL  FILL_4162
timestamp 1714281807
transform 1 0 1728 0 -1 170
box -8 -3 16 105
use FILL  FILL_4163
timestamp 1714281807
transform 1 0 1720 0 -1 170
box -8 -3 16 105
use FILL  FILL_4164
timestamp 1714281807
transform 1 0 1712 0 -1 170
box -8 -3 16 105
use FILL  FILL_4165
timestamp 1714281807
transform 1 0 1680 0 -1 170
box -8 -3 16 105
use FILL  FILL_4166
timestamp 1714281807
transform 1 0 1672 0 -1 170
box -8 -3 16 105
use FILL  FILL_4167
timestamp 1714281807
transform 1 0 1568 0 -1 170
box -8 -3 16 105
use FILL  FILL_4168
timestamp 1714281807
transform 1 0 1560 0 -1 170
box -8 -3 16 105
use FILL  FILL_4169
timestamp 1714281807
transform 1 0 1552 0 -1 170
box -8 -3 16 105
use FILL  FILL_4170
timestamp 1714281807
transform 1 0 1520 0 -1 170
box -8 -3 16 105
use FILL  FILL_4171
timestamp 1714281807
transform 1 0 1512 0 -1 170
box -8 -3 16 105
use FILL  FILL_4172
timestamp 1714281807
transform 1 0 1408 0 -1 170
box -8 -3 16 105
use FILL  FILL_4173
timestamp 1714281807
transform 1 0 1400 0 -1 170
box -8 -3 16 105
use FILL  FILL_4174
timestamp 1714281807
transform 1 0 1392 0 -1 170
box -8 -3 16 105
use FILL  FILL_4175
timestamp 1714281807
transform 1 0 1384 0 -1 170
box -8 -3 16 105
use FILL  FILL_4176
timestamp 1714281807
transform 1 0 1352 0 -1 170
box -8 -3 16 105
use FILL  FILL_4177
timestamp 1714281807
transform 1 0 1344 0 -1 170
box -8 -3 16 105
use FILL  FILL_4178
timestamp 1714281807
transform 1 0 1336 0 -1 170
box -8 -3 16 105
use FILL  FILL_4179
timestamp 1714281807
transform 1 0 1232 0 -1 170
box -8 -3 16 105
use FILL  FILL_4180
timestamp 1714281807
transform 1 0 1224 0 -1 170
box -8 -3 16 105
use FILL  FILL_4181
timestamp 1714281807
transform 1 0 1216 0 -1 170
box -8 -3 16 105
use FILL  FILL_4182
timestamp 1714281807
transform 1 0 1208 0 -1 170
box -8 -3 16 105
use FILL  FILL_4183
timestamp 1714281807
transform 1 0 1176 0 -1 170
box -8 -3 16 105
use FILL  FILL_4184
timestamp 1714281807
transform 1 0 1168 0 -1 170
box -8 -3 16 105
use FILL  FILL_4185
timestamp 1714281807
transform 1 0 1160 0 -1 170
box -8 -3 16 105
use FILL  FILL_4186
timestamp 1714281807
transform 1 0 1152 0 -1 170
box -8 -3 16 105
use FILL  FILL_4187
timestamp 1714281807
transform 1 0 1048 0 -1 170
box -8 -3 16 105
use FILL  FILL_4188
timestamp 1714281807
transform 1 0 1040 0 -1 170
box -8 -3 16 105
use FILL  FILL_4189
timestamp 1714281807
transform 1 0 936 0 -1 170
box -8 -3 16 105
use FILL  FILL_4190
timestamp 1714281807
transform 1 0 928 0 -1 170
box -8 -3 16 105
use FILL  FILL_4191
timestamp 1714281807
transform 1 0 920 0 -1 170
box -8 -3 16 105
use FILL  FILL_4192
timestamp 1714281807
transform 1 0 912 0 -1 170
box -8 -3 16 105
use FILL  FILL_4193
timestamp 1714281807
transform 1 0 904 0 -1 170
box -8 -3 16 105
use FILL  FILL_4194
timestamp 1714281807
transform 1 0 896 0 -1 170
box -8 -3 16 105
use FILL  FILL_4195
timestamp 1714281807
transform 1 0 856 0 -1 170
box -8 -3 16 105
use FILL  FILL_4196
timestamp 1714281807
transform 1 0 848 0 -1 170
box -8 -3 16 105
use FILL  FILL_4197
timestamp 1714281807
transform 1 0 840 0 -1 170
box -8 -3 16 105
use FILL  FILL_4198
timestamp 1714281807
transform 1 0 832 0 -1 170
box -8 -3 16 105
use FILL  FILL_4199
timestamp 1714281807
transform 1 0 792 0 -1 170
box -8 -3 16 105
use FILL  FILL_4200
timestamp 1714281807
transform 1 0 784 0 -1 170
box -8 -3 16 105
use FILL  FILL_4201
timestamp 1714281807
transform 1 0 776 0 -1 170
box -8 -3 16 105
use FILL  FILL_4202
timestamp 1714281807
transform 1 0 768 0 -1 170
box -8 -3 16 105
use FILL  FILL_4203
timestamp 1714281807
transform 1 0 760 0 -1 170
box -8 -3 16 105
use FILL  FILL_4204
timestamp 1714281807
transform 1 0 720 0 -1 170
box -8 -3 16 105
use FILL  FILL_4205
timestamp 1714281807
transform 1 0 712 0 -1 170
box -8 -3 16 105
use FILL  FILL_4206
timestamp 1714281807
transform 1 0 704 0 -1 170
box -8 -3 16 105
use FILL  FILL_4207
timestamp 1714281807
transform 1 0 696 0 -1 170
box -8 -3 16 105
use FILL  FILL_4208
timestamp 1714281807
transform 1 0 656 0 -1 170
box -8 -3 16 105
use FILL  FILL_4209
timestamp 1714281807
transform 1 0 648 0 -1 170
box -8 -3 16 105
use FILL  FILL_4210
timestamp 1714281807
transform 1 0 640 0 -1 170
box -8 -3 16 105
use FILL  FILL_4211
timestamp 1714281807
transform 1 0 632 0 -1 170
box -8 -3 16 105
use FILL  FILL_4212
timestamp 1714281807
transform 1 0 624 0 -1 170
box -8 -3 16 105
use FILL  FILL_4213
timestamp 1714281807
transform 1 0 592 0 -1 170
box -8 -3 16 105
use FILL  FILL_4214
timestamp 1714281807
transform 1 0 584 0 -1 170
box -8 -3 16 105
use FILL  FILL_4215
timestamp 1714281807
transform 1 0 576 0 -1 170
box -8 -3 16 105
use FILL  FILL_4216
timestamp 1714281807
transform 1 0 568 0 -1 170
box -8 -3 16 105
use FILL  FILL_4217
timestamp 1714281807
transform 1 0 544 0 -1 170
box -8 -3 16 105
use FILL  FILL_4218
timestamp 1714281807
transform 1 0 536 0 -1 170
box -8 -3 16 105
use FILL  FILL_4219
timestamp 1714281807
transform 1 0 528 0 -1 170
box -8 -3 16 105
use FILL  FILL_4220
timestamp 1714281807
transform 1 0 488 0 -1 170
box -8 -3 16 105
use FILL  FILL_4221
timestamp 1714281807
transform 1 0 480 0 -1 170
box -8 -3 16 105
use FILL  FILL_4222
timestamp 1714281807
transform 1 0 472 0 -1 170
box -8 -3 16 105
use FILL  FILL_4223
timestamp 1714281807
transform 1 0 464 0 -1 170
box -8 -3 16 105
use FILL  FILL_4224
timestamp 1714281807
transform 1 0 456 0 -1 170
box -8 -3 16 105
use FILL  FILL_4225
timestamp 1714281807
transform 1 0 448 0 -1 170
box -8 -3 16 105
use FILL  FILL_4226
timestamp 1714281807
transform 1 0 392 0 -1 170
box -8 -3 16 105
use FILL  FILL_4227
timestamp 1714281807
transform 1 0 384 0 -1 170
box -8 -3 16 105
use FILL  FILL_4228
timestamp 1714281807
transform 1 0 376 0 -1 170
box -8 -3 16 105
use FILL  FILL_4229
timestamp 1714281807
transform 1 0 368 0 -1 170
box -8 -3 16 105
use FILL  FILL_4230
timestamp 1714281807
transform 1 0 360 0 -1 170
box -8 -3 16 105
use FILL  FILL_4231
timestamp 1714281807
transform 1 0 352 0 -1 170
box -8 -3 16 105
use FILL  FILL_4232
timestamp 1714281807
transform 1 0 312 0 -1 170
box -8 -3 16 105
use FILL  FILL_4233
timestamp 1714281807
transform 1 0 304 0 -1 170
box -8 -3 16 105
use FILL  FILL_4234
timestamp 1714281807
transform 1 0 296 0 -1 170
box -8 -3 16 105
use FILL  FILL_4235
timestamp 1714281807
transform 1 0 288 0 -1 170
box -8 -3 16 105
use FILL  FILL_4236
timestamp 1714281807
transform 1 0 280 0 -1 170
box -8 -3 16 105
use FILL  FILL_4237
timestamp 1714281807
transform 1 0 248 0 -1 170
box -8 -3 16 105
use FILL  FILL_4238
timestamp 1714281807
transform 1 0 240 0 -1 170
box -8 -3 16 105
use FILL  FILL_4239
timestamp 1714281807
transform 1 0 232 0 -1 170
box -8 -3 16 105
use FILL  FILL_4240
timestamp 1714281807
transform 1 0 224 0 -1 170
box -8 -3 16 105
use FILL  FILL_4241
timestamp 1714281807
transform 1 0 216 0 -1 170
box -8 -3 16 105
use FILL  FILL_4242
timestamp 1714281807
transform 1 0 208 0 -1 170
box -8 -3 16 105
use FILL  FILL_4243
timestamp 1714281807
transform 1 0 200 0 -1 170
box -8 -3 16 105
use FILL  FILL_4244
timestamp 1714281807
transform 1 0 192 0 -1 170
box -8 -3 16 105
use FILL  FILL_4245
timestamp 1714281807
transform 1 0 184 0 -1 170
box -8 -3 16 105
use FILL  FILL_4246
timestamp 1714281807
transform 1 0 176 0 -1 170
box -8 -3 16 105
use FILL  FILL_4247
timestamp 1714281807
transform 1 0 168 0 -1 170
box -8 -3 16 105
use FILL  FILL_4248
timestamp 1714281807
transform 1 0 160 0 -1 170
box -8 -3 16 105
use FILL  FILL_4249
timestamp 1714281807
transform 1 0 152 0 -1 170
box -8 -3 16 105
use FILL  FILL_4250
timestamp 1714281807
transform 1 0 144 0 -1 170
box -8 -3 16 105
use FILL  FILL_4251
timestamp 1714281807
transform 1 0 136 0 -1 170
box -8 -3 16 105
use FILL  FILL_4252
timestamp 1714281807
transform 1 0 128 0 -1 170
box -8 -3 16 105
use FILL  FILL_4253
timestamp 1714281807
transform 1 0 120 0 -1 170
box -8 -3 16 105
use FILL  FILL_4254
timestamp 1714281807
transform 1 0 112 0 -1 170
box -8 -3 16 105
use FILL  FILL_4255
timestamp 1714281807
transform 1 0 104 0 -1 170
box -8 -3 16 105
use FILL  FILL_4256
timestamp 1714281807
transform 1 0 96 0 -1 170
box -8 -3 16 105
use FILL  FILL_4257
timestamp 1714281807
transform 1 0 88 0 -1 170
box -8 -3 16 105
use FILL  FILL_4258
timestamp 1714281807
transform 1 0 80 0 -1 170
box -8 -3 16 105
use FILL  FILL_4259
timestamp 1714281807
transform 1 0 72 0 -1 170
box -8 -3 16 105
use INVX2  INVX2_0
timestamp 1714281807
transform 1 0 584 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_1
timestamp 1714281807
transform 1 0 1184 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_2
timestamp 1714281807
transform 1 0 416 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_3
timestamp 1714281807
transform 1 0 416 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_4
timestamp 1714281807
transform 1 0 544 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_5
timestamp 1714281807
transform 1 0 1048 0 1 970
box -9 -3 26 105
use INVX2  INVX2_6
timestamp 1714281807
transform 1 0 1080 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_7
timestamp 1714281807
transform 1 0 432 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_8
timestamp 1714281807
transform 1 0 1240 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_9
timestamp 1714281807
transform 1 0 1160 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_10
timestamp 1714281807
transform 1 0 1024 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_11
timestamp 1714281807
transform 1 0 1224 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_12
timestamp 1714281807
transform 1 0 1064 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_13
timestamp 1714281807
transform 1 0 1192 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_14
timestamp 1714281807
transform 1 0 912 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_15
timestamp 1714281807
transform 1 0 992 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_16
timestamp 1714281807
transform 1 0 1144 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_17
timestamp 1714281807
transform 1 0 1200 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_18
timestamp 1714281807
transform 1 0 472 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_19
timestamp 1714281807
transform 1 0 288 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_20
timestamp 1714281807
transform 1 0 312 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_21
timestamp 1714281807
transform 1 0 464 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_22
timestamp 1714281807
transform 1 0 1056 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_23
timestamp 1714281807
transform 1 0 784 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_24
timestamp 1714281807
transform 1 0 664 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_25
timestamp 1714281807
transform 1 0 688 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_26
timestamp 1714281807
transform 1 0 888 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_27
timestamp 1714281807
transform 1 0 736 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_28
timestamp 1714281807
transform 1 0 584 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_29
timestamp 1714281807
transform 1 0 352 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_30
timestamp 1714281807
transform 1 0 296 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_31
timestamp 1714281807
transform 1 0 192 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_32
timestamp 1714281807
transform 1 0 240 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_33
timestamp 1714281807
transform 1 0 440 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_34
timestamp 1714281807
transform 1 0 624 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_35
timestamp 1714281807
transform 1 0 760 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_36
timestamp 1714281807
transform 1 0 1152 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_37
timestamp 1714281807
transform 1 0 1008 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_38
timestamp 1714281807
transform 1 0 456 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_39
timestamp 1714281807
transform 1 0 2744 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_40
timestamp 1714281807
transform 1 0 2768 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_41
timestamp 1714281807
transform 1 0 2792 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_42
timestamp 1714281807
transform 1 0 856 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_43
timestamp 1714281807
transform 1 0 1416 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_44
timestamp 1714281807
transform 1 0 1344 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_45
timestamp 1714281807
transform 1 0 1032 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_46
timestamp 1714281807
transform 1 0 1432 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_47
timestamp 1714281807
transform 1 0 1344 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_48
timestamp 1714281807
transform 1 0 840 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_49
timestamp 1714281807
transform 1 0 712 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_50
timestamp 1714281807
transform 1 0 1440 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_51
timestamp 1714281807
transform 1 0 936 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_52
timestamp 1714281807
transform 1 0 800 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_53
timestamp 1714281807
transform 1 0 192 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_54
timestamp 1714281807
transform 1 0 192 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_55
timestamp 1714281807
transform 1 0 336 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_56
timestamp 1714281807
transform 1 0 336 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_57
timestamp 1714281807
transform 1 0 272 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_58
timestamp 1714281807
transform 1 0 200 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_59
timestamp 1714281807
transform 1 0 304 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_60
timestamp 1714281807
transform 1 0 392 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_61
timestamp 1714281807
transform 1 0 528 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_62
timestamp 1714281807
transform 1 0 320 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_63
timestamp 1714281807
transform 1 0 2232 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_64
timestamp 1714281807
transform 1 0 2088 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_65
timestamp 1714281807
transform 1 0 2288 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_66
timestamp 1714281807
transform 1 0 2704 0 1 570
box -9 -3 26 105
use INVX2  INVX2_67
timestamp 1714281807
transform 1 0 2872 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_68
timestamp 1714281807
transform 1 0 2760 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_69
timestamp 1714281807
transform 1 0 2096 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_70
timestamp 1714281807
transform 1 0 2264 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_71
timestamp 1714281807
transform 1 0 2392 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_72
timestamp 1714281807
transform 1 0 2688 0 1 170
box -9 -3 26 105
use INVX2  INVX2_73
timestamp 1714281807
transform 1 0 2872 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_74
timestamp 1714281807
transform 1 0 2872 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_75
timestamp 1714281807
transform 1 0 2216 0 1 970
box -9 -3 26 105
use INVX2  INVX2_76
timestamp 1714281807
transform 1 0 2376 0 1 970
box -9 -3 26 105
use INVX2  INVX2_77
timestamp 1714281807
transform 1 0 2344 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_78
timestamp 1714281807
transform 1 0 2680 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_79
timestamp 1714281807
transform 1 0 2872 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_80
timestamp 1714281807
transform 1 0 2920 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_81
timestamp 1714281807
transform 1 0 1480 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_82
timestamp 1714281807
transform 1 0 1352 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_83
timestamp 1714281807
transform 1 0 1344 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_84
timestamp 1714281807
transform 1 0 1728 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_85
timestamp 1714281807
transform 1 0 1856 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_86
timestamp 1714281807
transform 1 0 1960 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_87
timestamp 1714281807
transform 1 0 2584 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_88
timestamp 1714281807
transform 1 0 2720 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_89
timestamp 1714281807
transform 1 0 2856 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_90
timestamp 1714281807
transform 1 0 1792 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_91
timestamp 1714281807
transform 1 0 1904 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_92
timestamp 1714281807
transform 1 0 2016 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_93
timestamp 1714281807
transform 1 0 2104 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_94
timestamp 1714281807
transform 1 0 2232 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_95
timestamp 1714281807
transform 1 0 2360 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_96
timestamp 1714281807
transform 1 0 2736 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_97
timestamp 1714281807
transform 1 0 2872 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_98
timestamp 1714281807
transform 1 0 2824 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_99
timestamp 1714281807
transform 1 0 2544 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_100
timestamp 1714281807
transform 1 0 2800 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_101
timestamp 1714281807
transform 1 0 2672 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_102
timestamp 1714281807
transform 1 0 2536 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_103
timestamp 1714281807
transform 1 0 2648 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_104
timestamp 1714281807
transform 1 0 2792 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_105
timestamp 1714281807
transform 1 0 2440 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_106
timestamp 1714281807
transform 1 0 2536 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_107
timestamp 1714281807
transform 1 0 2296 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_108
timestamp 1714281807
transform 1 0 1936 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_109
timestamp 1714281807
transform 1 0 2072 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_110
timestamp 1714281807
transform 1 0 2056 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_111
timestamp 1714281807
transform 1 0 2032 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_112
timestamp 1714281807
transform 1 0 1928 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_113
timestamp 1714281807
transform 1 0 1928 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_114
timestamp 1714281807
transform 1 0 1424 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_115
timestamp 1714281807
transform 1 0 1344 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_116
timestamp 1714281807
transform 1 0 1432 0 1 770
box -9 -3 26 105
use INVX2  INVX2_117
timestamp 1714281807
transform 1 0 1520 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_118
timestamp 1714281807
transform 1 0 1576 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_119
timestamp 1714281807
transform 1 0 1504 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_120
timestamp 1714281807
transform 1 0 1360 0 1 570
box -9 -3 26 105
use INVX2  INVX2_121
timestamp 1714281807
transform 1 0 1640 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_122
timestamp 1714281807
transform 1 0 1368 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_123
timestamp 1714281807
transform 1 0 1920 0 1 770
box -9 -3 26 105
use INVX2  INVX2_124
timestamp 1714281807
transform 1 0 1944 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_125
timestamp 1714281807
transform 1 0 1704 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_126
timestamp 1714281807
transform 1 0 1768 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_127
timestamp 1714281807
transform 1 0 2160 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_128
timestamp 1714281807
transform 1 0 2040 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_129
timestamp 1714281807
transform 1 0 2288 0 1 570
box -9 -3 26 105
use INVX2  INVX2_130
timestamp 1714281807
transform 1 0 2544 0 1 570
box -9 -3 26 105
use INVX2  INVX2_131
timestamp 1714281807
transform 1 0 2496 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_132
timestamp 1714281807
transform 1 0 2248 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_133
timestamp 1714281807
transform 1 0 2472 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_134
timestamp 1714281807
transform 1 0 2344 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_135
timestamp 1714281807
transform 1 0 1000 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_136
timestamp 1714281807
transform 1 0 472 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_137
timestamp 1714281807
transform 1 0 464 0 1 970
box -9 -3 26 105
use INVX2  INVX2_138
timestamp 1714281807
transform 1 0 720 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_139
timestamp 1714281807
transform 1 0 896 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_140
timestamp 1714281807
transform 1 0 936 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_141
timestamp 1714281807
transform 1 0 992 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_142
timestamp 1714281807
transform 1 0 1168 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_143
timestamp 1714281807
transform 1 0 1072 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_144
timestamp 1714281807
transform 1 0 448 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_145
timestamp 1714281807
transform 1 0 384 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_146
timestamp 1714281807
transform 1 0 1792 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_147
timestamp 1714281807
transform 1 0 1536 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_148
timestamp 1714281807
transform 1 0 1624 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_149
timestamp 1714281807
transform 1 0 1816 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_150
timestamp 1714281807
transform 1 0 1672 0 1 970
box -9 -3 26 105
use INVX2  INVX2_151
timestamp 1714281807
transform 1 0 1816 0 1 970
box -9 -3 26 105
use INVX2  INVX2_152
timestamp 1714281807
transform 1 0 1368 0 1 970
box -9 -3 26 105
use INVX2  INVX2_153
timestamp 1714281807
transform 1 0 1080 0 1 570
box -9 -3 26 105
use INVX2  INVX2_154
timestamp 1714281807
transform 1 0 1064 0 1 770
box -9 -3 26 105
use INVX2  INVX2_155
timestamp 1714281807
transform 1 0 1208 0 1 170
box -9 -3 26 105
use INVX2  INVX2_156
timestamp 1714281807
transform 1 0 1168 0 1 170
box -9 -3 26 105
use INVX2  INVX2_157
timestamp 1714281807
transform 1 0 1024 0 1 370
box -9 -3 26 105
use INVX2  INVX2_158
timestamp 1714281807
transform 1 0 1360 0 1 170
box -9 -3 26 105
use INVX2  INVX2_159
timestamp 1714281807
transform 1 0 1752 0 1 170
box -9 -3 26 105
use INVX2  INVX2_160
timestamp 1714281807
transform 1 0 1504 0 1 170
box -9 -3 26 105
use INVX2  INVX2_161
timestamp 1714281807
transform 1 0 1808 0 1 170
box -9 -3 26 105
use INVX2  INVX2_162
timestamp 1714281807
transform 1 0 2064 0 1 170
box -9 -3 26 105
use INVX2  INVX2_163
timestamp 1714281807
transform 1 0 2088 0 1 170
box -9 -3 26 105
use INVX2  INVX2_164
timestamp 1714281807
transform 1 0 2240 0 1 170
box -9 -3 26 105
use INVX2  INVX2_165
timestamp 1714281807
transform 1 0 2624 0 1 170
box -9 -3 26 105
use INVX2  INVX2_166
timestamp 1714281807
transform 1 0 2408 0 1 170
box -9 -3 26 105
use INVX2  INVX2_167
timestamp 1714281807
transform 1 0 1944 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_168
timestamp 1714281807
transform 1 0 1872 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_169
timestamp 1714281807
transform 1 0 1656 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_170
timestamp 1714281807
transform 1 0 536 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_171
timestamp 1714281807
transform 1 0 1416 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_172
timestamp 1714281807
transform 1 0 648 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_173
timestamp 1714281807
transform 1 0 696 0 1 970
box -9 -3 26 105
use INVX2  INVX2_174
timestamp 1714281807
transform 1 0 768 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_175
timestamp 1714281807
transform 1 0 1856 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_176
timestamp 1714281807
transform 1 0 1624 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_177
timestamp 1714281807
transform 1 0 2024 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_178
timestamp 1714281807
transform 1 0 1896 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_179
timestamp 1714281807
transform 1 0 1712 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_180
timestamp 1714281807
transform 1 0 1736 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_181
timestamp 1714281807
transform 1 0 1704 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_182
timestamp 1714281807
transform 1 0 616 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_183
timestamp 1714281807
transform 1 0 472 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_184
timestamp 1714281807
transform 1 0 1032 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_185
timestamp 1714281807
transform 1 0 1000 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_186
timestamp 1714281807
transform 1 0 656 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_187
timestamp 1714281807
transform 1 0 624 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_188
timestamp 1714281807
transform 1 0 760 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_189
timestamp 1714281807
transform 1 0 752 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_190
timestamp 1714281807
transform 1 0 560 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_191
timestamp 1714281807
transform 1 0 744 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_192
timestamp 1714281807
transform 1 0 776 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_193
timestamp 1714281807
transform 1 0 600 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_194
timestamp 1714281807
transform 1 0 1192 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_195
timestamp 1714281807
transform 1 0 1232 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_196
timestamp 1714281807
transform 1 0 1144 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_197
timestamp 1714281807
transform 1 0 1344 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_198
timestamp 1714281807
transform 1 0 1224 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_199
timestamp 1714281807
transform 1 0 1096 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_200
timestamp 1714281807
transform 1 0 1296 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_201
timestamp 1714281807
transform 1 0 1200 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_202
timestamp 1714281807
transform 1 0 912 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_203
timestamp 1714281807
transform 1 0 792 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_204
timestamp 1714281807
transform 1 0 896 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_205
timestamp 1714281807
transform 1 0 992 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_206
timestamp 1714281807
transform 1 0 856 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_207
timestamp 1714281807
transform 1 0 960 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_208
timestamp 1714281807
transform 1 0 664 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_209
timestamp 1714281807
transform 1 0 856 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_210
timestamp 1714281807
transform 1 0 776 0 1 970
box -9 -3 26 105
use INVX2  INVX2_211
timestamp 1714281807
transform 1 0 272 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_212
timestamp 1714281807
transform 1 0 688 0 1 570
box -9 -3 26 105
use INVX2  INVX2_213
timestamp 1714281807
transform 1 0 792 0 1 570
box -9 -3 26 105
use INVX2  INVX2_214
timestamp 1714281807
transform 1 0 352 0 1 370
box -9 -3 26 105
use INVX2  INVX2_215
timestamp 1714281807
transform 1 0 424 0 1 170
box -9 -3 26 105
use INVX2  INVX2_216
timestamp 1714281807
transform 1 0 400 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_217
timestamp 1714281807
transform 1 0 672 0 1 170
box -9 -3 26 105
use INVX2  INVX2_218
timestamp 1714281807
transform 1 0 640 0 1 170
box -9 -3 26 105
use INVX2  INVX2_219
timestamp 1714281807
transform 1 0 544 0 1 370
box -9 -3 26 105
use INVX2  INVX2_220
timestamp 1714281807
transform 1 0 552 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_221
timestamp 1714281807
transform 1 0 376 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_222
timestamp 1714281807
transform 1 0 872 0 -1 370
box -9 -3 26 105
use M2_M1  M2_M1_0
timestamp 1714281807
transform 1 0 1148 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1
timestamp 1714281807
transform 1 0 948 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2
timestamp 1714281807
transform 1 0 860 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3
timestamp 1714281807
transform 1 0 836 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_4
timestamp 1714281807
transform 1 0 732 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5
timestamp 1714281807
transform 1 0 700 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6
timestamp 1714281807
transform 1 0 636 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_7
timestamp 1714281807
transform 1 0 628 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_8
timestamp 1714281807
transform 1 0 500 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_9
timestamp 1714281807
transform 1 0 436 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_10
timestamp 1714281807
transform 1 0 412 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_11
timestamp 1714281807
transform 1 0 412 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_12
timestamp 1714281807
transform 1 0 604 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_13
timestamp 1714281807
transform 1 0 588 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_14
timestamp 1714281807
transform 1 0 532 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_15
timestamp 1714281807
transform 1 0 780 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_16
timestamp 1714281807
transform 1 0 740 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_17
timestamp 1714281807
transform 1 0 932 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_18
timestamp 1714281807
transform 1 0 892 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_19
timestamp 1714281807
transform 1 0 1308 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_20
timestamp 1714281807
transform 1 0 1204 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_21
timestamp 1714281807
transform 1 0 1252 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_22
timestamp 1714281807
transform 1 0 1148 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_23
timestamp 1714281807
transform 1 0 1100 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_24
timestamp 1714281807
transform 1 0 996 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_25
timestamp 1714281807
transform 1 0 468 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_26
timestamp 1714281807
transform 1 0 412 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_27
timestamp 1714281807
transform 1 0 316 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_28
timestamp 1714281807
transform 1 0 276 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_29
timestamp 1714281807
transform 1 0 2124 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_30
timestamp 1714281807
transform 1 0 2052 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_31
timestamp 1714281807
transform 1 0 1668 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_32
timestamp 1714281807
transform 1 0 1652 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_33
timestamp 1714281807
transform 1 0 2052 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_34
timestamp 1714281807
transform 1 0 2052 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_35
timestamp 1714281807
transform 1 0 1724 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_36
timestamp 1714281807
transform 1 0 1620 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_37
timestamp 1714281807
transform 1 0 1996 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_38
timestamp 1714281807
transform 1 0 1900 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_39
timestamp 1714281807
transform 1 0 1852 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_40
timestamp 1714281807
transform 1 0 1740 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_41
timestamp 1714281807
transform 1 0 1972 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_42
timestamp 1714281807
transform 1 0 1860 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_43
timestamp 1714281807
transform 1 0 1812 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_44
timestamp 1714281807
transform 1 0 1812 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_45
timestamp 1714281807
transform 1 0 2028 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_46
timestamp 1714281807
transform 1 0 1932 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_47
timestamp 1714281807
transform 1 0 1652 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_48
timestamp 1714281807
transform 1 0 1652 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_49
timestamp 1714281807
transform 1 0 2036 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_50
timestamp 1714281807
transform 1 0 1980 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_51
timestamp 1714281807
transform 1 0 1772 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_52
timestamp 1714281807
transform 1 0 1412 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_53
timestamp 1714281807
transform 1 0 1412 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_54
timestamp 1714281807
transform 1 0 1292 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_55
timestamp 1714281807
transform 1 0 1180 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_56
timestamp 1714281807
transform 1 0 1332 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_57
timestamp 1714281807
transform 1 0 1164 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_58
timestamp 1714281807
transform 1 0 1156 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_59
timestamp 1714281807
transform 1 0 1508 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_60
timestamp 1714281807
transform 1 0 1420 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_61
timestamp 1714281807
transform 1 0 1236 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_62
timestamp 1714281807
transform 1 0 1348 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_63
timestamp 1714281807
transform 1 0 1180 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_64
timestamp 1714281807
transform 1 0 1140 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_65
timestamp 1714281807
transform 1 0 1676 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_66
timestamp 1714281807
transform 1 0 1644 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_67
timestamp 1714281807
transform 1 0 1372 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_68
timestamp 1714281807
transform 1 0 1188 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_69
timestamp 1714281807
transform 1 0 1340 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_70
timestamp 1714281807
transform 1 0 1276 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_71
timestamp 1714281807
transform 1 0 1252 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_72
timestamp 1714281807
transform 1 0 1820 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_73
timestamp 1714281807
transform 1 0 1700 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_74
timestamp 1714281807
transform 1 0 1588 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_75
timestamp 1714281807
transform 1 0 1540 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_76
timestamp 1714281807
transform 1 0 1980 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_77
timestamp 1714281807
transform 1 0 1924 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_78
timestamp 1714281807
transform 1 0 1780 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_79
timestamp 1714281807
transform 1 0 1692 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_80
timestamp 1714281807
transform 1 0 1900 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_81
timestamp 1714281807
transform 1 0 1892 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_82
timestamp 1714281807
transform 1 0 1420 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_83
timestamp 1714281807
transform 1 0 2756 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_84
timestamp 1714281807
transform 1 0 2740 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_85
timestamp 1714281807
transform 1 0 2924 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_86
timestamp 1714281807
transform 1 0 2868 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_87
timestamp 1714281807
transform 1 0 2852 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_88
timestamp 1714281807
transform 1 0 2812 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_89
timestamp 1714281807
transform 1 0 2756 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_90
timestamp 1714281807
transform 1 0 2716 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_91
timestamp 1714281807
transform 1 0 2708 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_92
timestamp 1714281807
transform 1 0 2700 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_93
timestamp 1714281807
transform 1 0 2700 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_94
timestamp 1714281807
transform 1 0 2036 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_95
timestamp 1714281807
transform 1 0 2028 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_96
timestamp 1714281807
transform 1 0 2012 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_97
timestamp 1714281807
transform 1 0 2004 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_98
timestamp 1714281807
transform 1 0 2228 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_99
timestamp 1714281807
transform 1 0 2204 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_100
timestamp 1714281807
transform 1 0 2124 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_101
timestamp 1714281807
transform 1 0 2092 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_102
timestamp 1714281807
transform 1 0 1892 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_103
timestamp 1714281807
transform 1 0 1844 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_104
timestamp 1714281807
transform 1 0 1836 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_105
timestamp 1714281807
transform 1 0 1772 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_106
timestamp 1714281807
transform 1 0 2468 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_107
timestamp 1714281807
transform 1 0 2460 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_108
timestamp 1714281807
transform 1 0 2460 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_109
timestamp 1714281807
transform 1 0 2644 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_110
timestamp 1714281807
transform 1 0 2548 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_111
timestamp 1714281807
transform 1 0 2540 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_112
timestamp 1714281807
transform 1 0 2540 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_113
timestamp 1714281807
transform 1 0 2356 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_114
timestamp 1714281807
transform 1 0 2268 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_115
timestamp 1714281807
transform 1 0 2268 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_116
timestamp 1714281807
transform 1 0 2260 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_117
timestamp 1714281807
transform 1 0 2476 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_118
timestamp 1714281807
transform 1 0 2412 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_119
timestamp 1714281807
transform 1 0 2292 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_120
timestamp 1714281807
transform 1 0 2292 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_121
timestamp 1714281807
transform 1 0 2484 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_122
timestamp 1714281807
transform 1 0 2476 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_123
timestamp 1714281807
transform 1 0 2436 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_124
timestamp 1714281807
transform 1 0 2292 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_125
timestamp 1714281807
transform 1 0 2436 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_126
timestamp 1714281807
transform 1 0 2428 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_127
timestamp 1714281807
transform 1 0 2220 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_128
timestamp 1714281807
transform 1 0 2180 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_129
timestamp 1714281807
transform 1 0 2900 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_130
timestamp 1714281807
transform 1 0 2796 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_131
timestamp 1714281807
transform 1 0 2796 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_132
timestamp 1714281807
transform 1 0 2684 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_133
timestamp 1714281807
transform 1 0 2660 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_134
timestamp 1714281807
transform 1 0 2660 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_135
timestamp 1714281807
transform 1 0 2652 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_136
timestamp 1714281807
transform 1 0 2620 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_137
timestamp 1714281807
transform 1 0 2524 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_138
timestamp 1714281807
transform 1 0 2516 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_139
timestamp 1714281807
transform 1 0 2900 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_140
timestamp 1714281807
transform 1 0 2748 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_141
timestamp 1714281807
transform 1 0 2692 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_142
timestamp 1714281807
transform 1 0 2676 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_143
timestamp 1714281807
transform 1 0 2844 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_144
timestamp 1714281807
transform 1 0 2804 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_145
timestamp 1714281807
transform 1 0 2780 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_146
timestamp 1714281807
transform 1 0 2772 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_147
timestamp 1714281807
transform 1 0 2748 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_148
timestamp 1714281807
transform 1 0 2724 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_149
timestamp 1714281807
transform 1 0 2580 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_150
timestamp 1714281807
transform 1 0 2548 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_151
timestamp 1714281807
transform 1 0 2548 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_152
timestamp 1714281807
transform 1 0 1556 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_153
timestamp 1714281807
transform 1 0 1492 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_154
timestamp 1714281807
transform 1 0 1484 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_155
timestamp 1714281807
transform 1 0 1396 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_156
timestamp 1714281807
transform 1 0 1628 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_157
timestamp 1714281807
transform 1 0 1580 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_158
timestamp 1714281807
transform 1 0 1524 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_159
timestamp 1714281807
transform 1 0 1420 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_160
timestamp 1714281807
transform 1 0 1564 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_161
timestamp 1714281807
transform 1 0 1548 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_162
timestamp 1714281807
transform 1 0 1524 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_163
timestamp 1714281807
transform 1 0 1468 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_164
timestamp 1714281807
transform 1 0 2020 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_165
timestamp 1714281807
transform 1 0 1940 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_166
timestamp 1714281807
transform 1 0 1924 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_167
timestamp 1714281807
transform 1 0 1924 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_168
timestamp 1714281807
transform 1 0 1908 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_169
timestamp 1714281807
transform 1 0 1844 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_170
timestamp 1714281807
transform 1 0 1804 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_171
timestamp 1714281807
transform 1 0 1852 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_172
timestamp 1714281807
transform 1 0 1836 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_173
timestamp 1714281807
transform 1 0 1724 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_174
timestamp 1714281807
transform 1 0 1724 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_175
timestamp 1714281807
transform 1 0 2388 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_176
timestamp 1714281807
transform 1 0 2380 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_177
timestamp 1714281807
transform 1 0 2380 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_178
timestamp 1714281807
transform 1 0 2276 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_179
timestamp 1714281807
transform 1 0 2276 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_180
timestamp 1714281807
transform 1 0 2268 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_181
timestamp 1714281807
transform 1 0 2164 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_182
timestamp 1714281807
transform 1 0 2164 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_183
timestamp 1714281807
transform 1 0 2060 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_184
timestamp 1714281807
transform 1 0 2060 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_185
timestamp 1714281807
transform 1 0 2796 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_186
timestamp 1714281807
transform 1 0 2772 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_187
timestamp 1714281807
transform 1 0 2708 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_188
timestamp 1714281807
transform 1 0 2708 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_189
timestamp 1714281807
transform 1 0 2764 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_190
timestamp 1714281807
transform 1 0 2724 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_191
timestamp 1714281807
transform 1 0 2700 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_192
timestamp 1714281807
transform 1 0 2676 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_193
timestamp 1714281807
transform 1 0 2740 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_194
timestamp 1714281807
transform 1 0 2724 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_195
timestamp 1714281807
transform 1 0 2724 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_196
timestamp 1714281807
transform 1 0 2708 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_197
timestamp 1714281807
transform 1 0 2484 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_198
timestamp 1714281807
transform 1 0 2292 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_199
timestamp 1714281807
transform 1 0 2292 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_200
timestamp 1714281807
transform 1 0 2292 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_201
timestamp 1714281807
transform 1 0 2356 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_202
timestamp 1714281807
transform 1 0 2204 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_203
timestamp 1714281807
transform 1 0 2092 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_204
timestamp 1714281807
transform 1 0 2380 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_205
timestamp 1714281807
transform 1 0 2300 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_206
timestamp 1714281807
transform 1 0 2284 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_207
timestamp 1714281807
transform 1 0 2236 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_208
timestamp 1714281807
transform 1 0 404 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_209
timestamp 1714281807
transform 1 0 388 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_210
timestamp 1714281807
transform 1 0 388 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_211
timestamp 1714281807
transform 1 0 388 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_212
timestamp 1714281807
transform 1 0 516 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_213
timestamp 1714281807
transform 1 0 452 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_214
timestamp 1714281807
transform 1 0 452 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_215
timestamp 1714281807
transform 1 0 996 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_216
timestamp 1714281807
transform 1 0 988 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_217
timestamp 1714281807
transform 1 0 980 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_218
timestamp 1714281807
transform 1 0 964 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_219
timestamp 1714281807
transform 1 0 892 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_220
timestamp 1714281807
transform 1 0 628 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_221
timestamp 1714281807
transform 1 0 620 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_222
timestamp 1714281807
transform 1 0 876 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_223
timestamp 1714281807
transform 1 0 860 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_224
timestamp 1714281807
transform 1 0 860 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_225
timestamp 1714281807
transform 1 0 812 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_226
timestamp 1714281807
transform 1 0 724 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_227
timestamp 1714281807
transform 1 0 1604 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_228
timestamp 1714281807
transform 1 0 1540 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_229
timestamp 1714281807
transform 1 0 1892 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_230
timestamp 1714281807
transform 1 0 1788 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_231
timestamp 1714281807
transform 1 0 1788 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_232
timestamp 1714281807
transform 1 0 1932 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_233
timestamp 1714281807
transform 1 0 1820 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_234
timestamp 1714281807
transform 1 0 1956 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_235
timestamp 1714281807
transform 1 0 1812 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_236
timestamp 1714281807
transform 1 0 1676 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_237
timestamp 1714281807
transform 1 0 1044 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_238
timestamp 1714281807
transform 1 0 1028 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_239
timestamp 1714281807
transform 1 0 1332 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_240
timestamp 1714281807
transform 1 0 1212 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_241
timestamp 1714281807
transform 1 0 1612 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_242
timestamp 1714281807
transform 1 0 1508 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_243
timestamp 1714281807
transform 1 0 1476 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_244
timestamp 1714281807
transform 1 0 1364 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_245
timestamp 1714281807
transform 1 0 2212 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_246
timestamp 1714281807
transform 1 0 2092 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_247
timestamp 1714281807
transform 1 0 1932 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_248
timestamp 1714281807
transform 1 0 1812 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_249
timestamp 1714281807
transform 1 0 2524 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_250
timestamp 1714281807
transform 1 0 2404 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_251
timestamp 1714281807
transform 1 0 2356 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_252
timestamp 1714281807
transform 1 0 2236 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_253
timestamp 1714281807
transform 1 0 2996 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_254
timestamp 1714281807
transform 1 0 2876 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_255
timestamp 1714281807
transform 1 0 2996 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_256
timestamp 1714281807
transform 1 0 2876 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_257
timestamp 1714281807
transform 1 0 2804 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_258
timestamp 1714281807
transform 1 0 2692 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_259
timestamp 1714281807
transform 1 0 2348 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_260
timestamp 1714281807
transform 1 0 2308 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_261
timestamp 1714281807
transform 1 0 2980 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_262
timestamp 1714281807
transform 1 0 2924 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_263
timestamp 1714281807
transform 1 0 2996 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_264
timestamp 1714281807
transform 1 0 2876 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_265
timestamp 1714281807
transform 1 0 1372 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_266
timestamp 1714281807
transform 1 0 1348 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_267
timestamp 1714281807
transform 1 0 2972 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_268
timestamp 1714281807
transform 1 0 2860 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_269
timestamp 1714281807
transform 1 0 2844 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_270
timestamp 1714281807
transform 1 0 2724 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_271
timestamp 1714281807
transform 1 0 2468 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_272
timestamp 1714281807
transform 1 0 2364 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_273
timestamp 1714281807
transform 1 0 2340 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_274
timestamp 1714281807
transform 1 0 2236 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_275
timestamp 1714281807
transform 1 0 2212 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_276
timestamp 1714281807
transform 1 0 2108 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_277
timestamp 1714281807
transform 1 0 2956 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_278
timestamp 1714281807
transform 1 0 2828 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_279
timestamp 1714281807
transform 1 0 2996 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_280
timestamp 1714281807
transform 1 0 2876 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_281
timestamp 1714281807
transform 1 0 2860 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_282
timestamp 1714281807
transform 1 0 2732 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_283
timestamp 1714281807
transform 1 0 2428 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_284
timestamp 1714281807
transform 1 0 2300 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_285
timestamp 1714281807
transform 1 0 2500 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_286
timestamp 1714281807
transform 1 0 2444 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_287
timestamp 1714281807
transform 1 0 636 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_288
timestamp 1714281807
transform 1 0 636 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_289
timestamp 1714281807
transform 1 0 580 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_290
timestamp 1714281807
transform 1 0 508 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_291
timestamp 1714281807
transform 1 0 484 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_292
timestamp 1714281807
transform 1 0 436 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_293
timestamp 1714281807
transform 1 0 476 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_294
timestamp 1714281807
transform 1 0 468 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_295
timestamp 1714281807
transform 1 0 332 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_296
timestamp 1714281807
transform 1 0 380 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_297
timestamp 1714281807
transform 1 0 252 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_298
timestamp 1714281807
transform 1 0 252 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_299
timestamp 1714281807
transform 1 0 228 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_300
timestamp 1714281807
transform 1 0 284 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_301
timestamp 1714281807
transform 1 0 236 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_302
timestamp 1714281807
transform 1 0 356 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_303
timestamp 1714281807
transform 1 0 340 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_304
timestamp 1714281807
transform 1 0 284 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_305
timestamp 1714281807
transform 1 0 260 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_306
timestamp 1714281807
transform 1 0 588 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_307
timestamp 1714281807
transform 1 0 500 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_308
timestamp 1714281807
transform 1 0 500 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_309
timestamp 1714281807
transform 1 0 892 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_310
timestamp 1714281807
transform 1 0 812 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_311
timestamp 1714281807
transform 1 0 1380 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_312
timestamp 1714281807
transform 1 0 924 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_313
timestamp 1714281807
transform 1 0 884 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_314
timestamp 1714281807
transform 1 0 780 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_315
timestamp 1714281807
transform 1 0 668 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_316
timestamp 1714281807
transform 1 0 916 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_317
timestamp 1714281807
transform 1 0 812 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_318
timestamp 1714281807
transform 1 0 804 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_319
timestamp 1714281807
transform 1 0 1388 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_320
timestamp 1714281807
transform 1 0 1212 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_321
timestamp 1714281807
transform 1 0 1100 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_322
timestamp 1714281807
transform 1 0 1180 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_323
timestamp 1714281807
transform 1 0 1116 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_324
timestamp 1714281807
transform 1 0 1204 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_325
timestamp 1714281807
transform 1 0 1148 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_326
timestamp 1714281807
transform 1 0 1012 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_327
timestamp 1714281807
transform 1 0 1180 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_328
timestamp 1714281807
transform 1 0 1108 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_329
timestamp 1714281807
transform 1 0 932 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_330
timestamp 1714281807
transform 1 0 876 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_331
timestamp 1714281807
transform 1 0 852 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_332
timestamp 1714281807
transform 1 0 852 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_333
timestamp 1714281807
transform 1 0 796 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_334
timestamp 1714281807
transform 1 0 660 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_335
timestamp 1714281807
transform 1 0 636 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_336
timestamp 1714281807
transform 1 0 724 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_337
timestamp 1714281807
transform 1 0 716 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_338
timestamp 1714281807
transform 1 0 716 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_339
timestamp 1714281807
transform 1 0 700 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_340
timestamp 1714281807
transform 1 0 652 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_341
timestamp 1714281807
transform 1 0 652 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_342
timestamp 1714281807
transform 1 0 620 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_343
timestamp 1714281807
transform 1 0 388 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_344
timestamp 1714281807
transform 1 0 292 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_345
timestamp 1714281807
transform 1 0 268 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_346
timestamp 1714281807
transform 1 0 252 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_347
timestamp 1714281807
transform 1 0 444 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_348
timestamp 1714281807
transform 1 0 292 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_349
timestamp 1714281807
transform 1 0 276 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_350
timestamp 1714281807
transform 1 0 276 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_351
timestamp 1714281807
transform 1 0 940 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_352
timestamp 1714281807
transform 1 0 836 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_353
timestamp 1714281807
transform 1 0 740 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_354
timestamp 1714281807
transform 1 0 644 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_355
timestamp 1714281807
transform 1 0 548 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_356
timestamp 1714281807
transform 1 0 452 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_357
timestamp 1714281807
transform 1 0 356 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_358
timestamp 1714281807
transform 1 0 964 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_359
timestamp 1714281807
transform 1 0 860 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_360
timestamp 1714281807
transform 1 0 804 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_361
timestamp 1714281807
transform 1 0 700 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_362
timestamp 1714281807
transform 1 0 276 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_363
timestamp 1714281807
transform 1 0 252 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_364
timestamp 1714281807
transform 1 0 244 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_365
timestamp 1714281807
transform 1 0 244 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_366
timestamp 1714281807
transform 1 0 236 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_367
timestamp 1714281807
transform 1 0 228 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_368
timestamp 1714281807
transform 1 0 212 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_369
timestamp 1714281807
transform 1 0 164 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_370
timestamp 1714281807
transform 1 0 132 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_371
timestamp 1714281807
transform 1 0 100 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_372
timestamp 1714281807
transform 1 0 2524 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_373
timestamp 1714281807
transform 1 0 2508 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_374
timestamp 1714281807
transform 1 0 2492 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_375
timestamp 1714281807
transform 1 0 2492 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_376
timestamp 1714281807
transform 1 0 2484 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_377
timestamp 1714281807
transform 1 0 2116 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_378
timestamp 1714281807
transform 1 0 1468 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_379
timestamp 1714281807
transform 1 0 1428 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_380
timestamp 1714281807
transform 1 0 1396 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_381
timestamp 1714281807
transform 1 0 1396 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_382
timestamp 1714281807
transform 1 0 1388 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_383
timestamp 1714281807
transform 1 0 748 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_384
timestamp 1714281807
transform 1 0 724 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_385
timestamp 1714281807
transform 1 0 716 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_386
timestamp 1714281807
transform 1 0 2788 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_387
timestamp 1714281807
transform 1 0 2684 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_388
timestamp 1714281807
transform 1 0 2580 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_389
timestamp 1714281807
transform 1 0 2580 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_390
timestamp 1714281807
transform 1 0 2476 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_391
timestamp 1714281807
transform 1 0 2308 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_392
timestamp 1714281807
transform 1 0 2228 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_393
timestamp 1714281807
transform 1 0 2140 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_394
timestamp 1714281807
transform 1 0 1988 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_395
timestamp 1714281807
transform 1 0 1892 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_396
timestamp 1714281807
transform 1 0 1676 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_397
timestamp 1714281807
transform 1 0 1660 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_398
timestamp 1714281807
transform 1 0 1612 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_399
timestamp 1714281807
transform 1 0 1580 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_400
timestamp 1714281807
transform 1 0 2916 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_401
timestamp 1714281807
transform 1 0 2916 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_402
timestamp 1714281807
transform 1 0 2836 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_403
timestamp 1714281807
transform 1 0 2764 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_404
timestamp 1714281807
transform 1 0 2732 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_405
timestamp 1714281807
transform 1 0 2628 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_406
timestamp 1714281807
transform 1 0 2628 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_407
timestamp 1714281807
transform 1 0 2596 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_408
timestamp 1714281807
transform 1 0 2500 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_409
timestamp 1714281807
transform 1 0 2484 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_410
timestamp 1714281807
transform 1 0 2484 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_411
timestamp 1714281807
transform 1 0 2308 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_412
timestamp 1714281807
transform 1 0 2132 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_413
timestamp 1714281807
transform 1 0 2108 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_414
timestamp 1714281807
transform 1 0 1900 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_415
timestamp 1714281807
transform 1 0 1748 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_416
timestamp 1714281807
transform 1 0 1748 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_417
timestamp 1714281807
transform 1 0 1740 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_418
timestamp 1714281807
transform 1 0 1636 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_419
timestamp 1714281807
transform 1 0 1588 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_420
timestamp 1714281807
transform 1 0 1428 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_421
timestamp 1714281807
transform 1 0 1252 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_422
timestamp 1714281807
transform 1 0 1076 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_423
timestamp 1714281807
transform 1 0 1068 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_424
timestamp 1714281807
transform 1 0 956 0 1 255
box -2 -2 2 2
use M2_M1  M2_M1_425
timestamp 1714281807
transform 1 0 956 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_426
timestamp 1714281807
transform 1 0 924 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_427
timestamp 1714281807
transform 1 0 924 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_428
timestamp 1714281807
transform 1 0 924 0 1 255
box -2 -2 2 2
use M2_M1  M2_M1_429
timestamp 1714281807
transform 1 0 916 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_430
timestamp 1714281807
transform 1 0 2884 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_431
timestamp 1714281807
transform 1 0 2876 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_432
timestamp 1714281807
transform 1 0 2876 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_433
timestamp 1714281807
transform 1 0 2356 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_434
timestamp 1714281807
transform 1 0 2244 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_435
timestamp 1714281807
transform 1 0 2156 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_436
timestamp 1714281807
transform 1 0 2132 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_437
timestamp 1714281807
transform 1 0 2084 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_438
timestamp 1714281807
transform 1 0 1996 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_439
timestamp 1714281807
transform 1 0 1756 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_440
timestamp 1714281807
transform 1 0 1748 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_441
timestamp 1714281807
transform 1 0 1724 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_442
timestamp 1714281807
transform 1 0 1620 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_443
timestamp 1714281807
transform 1 0 1588 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_444
timestamp 1714281807
transform 1 0 2884 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_445
timestamp 1714281807
transform 1 0 2884 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_446
timestamp 1714281807
transform 1 0 2828 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_447
timestamp 1714281807
transform 1 0 2788 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_448
timestamp 1714281807
transform 1 0 2540 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_449
timestamp 1714281807
transform 1 0 2476 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_450
timestamp 1714281807
transform 1 0 2292 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_451
timestamp 1714281807
transform 1 0 2004 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_452
timestamp 1714281807
transform 1 0 1988 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_453
timestamp 1714281807
transform 1 0 1756 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_454
timestamp 1714281807
transform 1 0 1740 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_455
timestamp 1714281807
transform 1 0 1660 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_456
timestamp 1714281807
transform 1 0 1628 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_457
timestamp 1714281807
transform 1 0 1620 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_458
timestamp 1714281807
transform 1 0 2868 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_459
timestamp 1714281807
transform 1 0 2860 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_460
timestamp 1714281807
transform 1 0 2788 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_461
timestamp 1714281807
transform 1 0 2588 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_462
timestamp 1714281807
transform 1 0 2580 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_463
timestamp 1714281807
transform 1 0 2548 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_464
timestamp 1714281807
transform 1 0 2356 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_465
timestamp 1714281807
transform 1 0 2188 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_466
timestamp 1714281807
transform 1 0 2172 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_467
timestamp 1714281807
transform 1 0 2124 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_468
timestamp 1714281807
transform 1 0 2084 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_469
timestamp 1714281807
transform 1 0 1836 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_470
timestamp 1714281807
transform 1 0 1580 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_471
timestamp 1714281807
transform 1 0 1572 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_472
timestamp 1714281807
transform 1 0 2180 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_473
timestamp 1714281807
transform 1 0 2180 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_474
timestamp 1714281807
transform 1 0 2092 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_475
timestamp 1714281807
transform 1 0 2076 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_476
timestamp 1714281807
transform 1 0 2036 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_477
timestamp 1714281807
transform 1 0 2020 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_478
timestamp 1714281807
transform 1 0 1868 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_479
timestamp 1714281807
transform 1 0 1668 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_480
timestamp 1714281807
transform 1 0 1548 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_481
timestamp 1714281807
transform 1 0 1532 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_482
timestamp 1714281807
transform 1 0 1532 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_483
timestamp 1714281807
transform 1 0 1524 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_484
timestamp 1714281807
transform 1 0 1524 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_485
timestamp 1714281807
transform 1 0 1476 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_486
timestamp 1714281807
transform 1 0 1412 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_487
timestamp 1714281807
transform 1 0 1308 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_488
timestamp 1714281807
transform 1 0 1300 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_489
timestamp 1714281807
transform 1 0 1212 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_490
timestamp 1714281807
transform 1 0 1188 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_491
timestamp 1714281807
transform 1 0 1116 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_492
timestamp 1714281807
transform 1 0 1076 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_493
timestamp 1714281807
transform 1 0 972 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_494
timestamp 1714281807
transform 1 0 932 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_495
timestamp 1714281807
transform 1 0 836 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_496
timestamp 1714281807
transform 1 0 620 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_497
timestamp 1714281807
transform 1 0 604 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_498
timestamp 1714281807
transform 1 0 516 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_499
timestamp 1714281807
transform 1 0 492 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_500
timestamp 1714281807
transform 1 0 1020 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_501
timestamp 1714281807
transform 1 0 948 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_502
timestamp 1714281807
transform 1 0 924 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_503
timestamp 1714281807
transform 1 0 2140 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_504
timestamp 1714281807
transform 1 0 2100 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_505
timestamp 1714281807
transform 1 0 2084 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_506
timestamp 1714281807
transform 1 0 2076 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_507
timestamp 1714281807
transform 1 0 1732 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_508
timestamp 1714281807
transform 1 0 1724 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_509
timestamp 1714281807
transform 1 0 1724 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_510
timestamp 1714281807
transform 1 0 1724 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_511
timestamp 1714281807
transform 1 0 1556 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_512
timestamp 1714281807
transform 1 0 1532 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_513
timestamp 1714281807
transform 1 0 1524 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_514
timestamp 1714281807
transform 1 0 1396 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_515
timestamp 1714281807
transform 1 0 436 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_516
timestamp 1714281807
transform 1 0 420 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_517
timestamp 1714281807
transform 1 0 420 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_518
timestamp 1714281807
transform 1 0 420 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_519
timestamp 1714281807
transform 1 0 396 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_520
timestamp 1714281807
transform 1 0 980 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_521
timestamp 1714281807
transform 1 0 940 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_522
timestamp 1714281807
transform 1 0 924 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_523
timestamp 1714281807
transform 1 0 916 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_524
timestamp 1714281807
transform 1 0 876 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_525
timestamp 1714281807
transform 1 0 796 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_526
timestamp 1714281807
transform 1 0 780 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_527
timestamp 1714281807
transform 1 0 740 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_528
timestamp 1714281807
transform 1 0 460 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_529
timestamp 1714281807
transform 1 0 460 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_530
timestamp 1714281807
transform 1 0 372 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_531
timestamp 1714281807
transform 1 0 356 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_532
timestamp 1714281807
transform 1 0 356 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_533
timestamp 1714281807
transform 1 0 1204 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_534
timestamp 1714281807
transform 1 0 1116 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_535
timestamp 1714281807
transform 1 0 1036 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_536
timestamp 1714281807
transform 1 0 1004 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_537
timestamp 1714281807
transform 1 0 884 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_538
timestamp 1714281807
transform 1 0 804 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_539
timestamp 1714281807
transform 1 0 740 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_540
timestamp 1714281807
transform 1 0 636 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_541
timestamp 1714281807
transform 1 0 540 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_542
timestamp 1714281807
transform 1 0 484 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_543
timestamp 1714281807
transform 1 0 484 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_544
timestamp 1714281807
transform 1 0 476 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_545
timestamp 1714281807
transform 1 0 436 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_546
timestamp 1714281807
transform 1 0 2460 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_547
timestamp 1714281807
transform 1 0 2452 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_548
timestamp 1714281807
transform 1 0 2372 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_549
timestamp 1714281807
transform 1 0 2340 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_550
timestamp 1714281807
transform 1 0 2324 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_551
timestamp 1714281807
transform 1 0 2268 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_552
timestamp 1714281807
transform 1 0 2148 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_553
timestamp 1714281807
transform 1 0 2068 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_554
timestamp 1714281807
transform 1 0 2028 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_555
timestamp 1714281807
transform 1 0 1972 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_556
timestamp 1714281807
transform 1 0 1844 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_557
timestamp 1714281807
transform 1 0 1772 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_558
timestamp 1714281807
transform 1 0 1764 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_559
timestamp 1714281807
transform 1 0 2036 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_560
timestamp 1714281807
transform 1 0 1996 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_561
timestamp 1714281807
transform 1 0 1996 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_562
timestamp 1714281807
transform 1 0 1972 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_563
timestamp 1714281807
transform 1 0 1684 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_564
timestamp 1714281807
transform 1 0 1540 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_565
timestamp 1714281807
transform 1 0 1516 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_566
timestamp 1714281807
transform 1 0 1508 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_567
timestamp 1714281807
transform 1 0 1444 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_568
timestamp 1714281807
transform 1 0 1428 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_569
timestamp 1714281807
transform 1 0 1420 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_570
timestamp 1714281807
transform 1 0 1412 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_571
timestamp 1714281807
transform 1 0 1412 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_572
timestamp 1714281807
transform 1 0 1388 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_573
timestamp 1714281807
transform 1 0 2668 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_574
timestamp 1714281807
transform 1 0 2652 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_575
timestamp 1714281807
transform 1 0 2564 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_576
timestamp 1714281807
transform 1 0 2548 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_577
timestamp 1714281807
transform 1 0 2500 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_578
timestamp 1714281807
transform 1 0 2476 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_579
timestamp 1714281807
transform 1 0 2132 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_580
timestamp 1714281807
transform 1 0 2132 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_581
timestamp 1714281807
transform 1 0 2092 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_582
timestamp 1714281807
transform 1 0 1988 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_583
timestamp 1714281807
transform 1 0 1956 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_584
timestamp 1714281807
transform 1 0 1884 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_585
timestamp 1714281807
transform 1 0 1788 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_586
timestamp 1714281807
transform 1 0 2756 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_587
timestamp 1714281807
transform 1 0 2748 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_588
timestamp 1714281807
transform 1 0 2740 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_589
timestamp 1714281807
transform 1 0 2716 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_590
timestamp 1714281807
transform 1 0 2716 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_591
timestamp 1714281807
transform 1 0 2708 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_592
timestamp 1714281807
transform 1 0 2684 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_593
timestamp 1714281807
transform 1 0 2356 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_594
timestamp 1714281807
transform 1 0 2292 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_595
timestamp 1714281807
transform 1 0 2196 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_596
timestamp 1714281807
transform 1 0 2188 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_597
timestamp 1714281807
transform 1 0 2148 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_598
timestamp 1714281807
transform 1 0 2140 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_599
timestamp 1714281807
transform 1 0 2140 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_600
timestamp 1714281807
transform 1 0 2124 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_601
timestamp 1714281807
transform 1 0 1036 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_602
timestamp 1714281807
transform 1 0 604 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_603
timestamp 1714281807
transform 1 0 604 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_604
timestamp 1714281807
transform 1 0 1084 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_605
timestamp 1714281807
transform 1 0 1028 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_606
timestamp 1714281807
transform 1 0 348 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_607
timestamp 1714281807
transform 1 0 332 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_608
timestamp 1714281807
transform 1 0 308 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_609
timestamp 1714281807
transform 1 0 308 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_610
timestamp 1714281807
transform 1 0 252 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_611
timestamp 1714281807
transform 1 0 1260 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_612
timestamp 1714281807
transform 1 0 1228 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_613
timestamp 1714281807
transform 1 0 828 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_614
timestamp 1714281807
transform 1 0 820 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_615
timestamp 1714281807
transform 1 0 700 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_616
timestamp 1714281807
transform 1 0 540 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_617
timestamp 1714281807
transform 1 0 540 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_618
timestamp 1714281807
transform 1 0 1292 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_619
timestamp 1714281807
transform 1 0 1292 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_620
timestamp 1714281807
transform 1 0 1284 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_621
timestamp 1714281807
transform 1 0 1252 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_622
timestamp 1714281807
transform 1 0 1228 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_623
timestamp 1714281807
transform 1 0 1220 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_624
timestamp 1714281807
transform 1 0 1500 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_625
timestamp 1714281807
transform 1 0 1492 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_626
timestamp 1714281807
transform 1 0 1492 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_627
timestamp 1714281807
transform 1 0 1484 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_628
timestamp 1714281807
transform 1 0 1436 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_629
timestamp 1714281807
transform 1 0 1420 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_630
timestamp 1714281807
transform 1 0 1412 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_631
timestamp 1714281807
transform 1 0 1404 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_632
timestamp 1714281807
transform 1 0 1380 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_633
timestamp 1714281807
transform 1 0 1380 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_634
timestamp 1714281807
transform 1 0 1364 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_635
timestamp 1714281807
transform 1 0 1340 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_636
timestamp 1714281807
transform 1 0 1340 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_637
timestamp 1714281807
transform 1 0 1308 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_638
timestamp 1714281807
transform 1 0 1284 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_639
timestamp 1714281807
transform 1 0 1540 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_640
timestamp 1714281807
transform 1 0 1500 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_641
timestamp 1714281807
transform 1 0 1476 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_642
timestamp 1714281807
transform 1 0 1364 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_643
timestamp 1714281807
transform 1 0 1124 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_644
timestamp 1714281807
transform 1 0 1124 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_645
timestamp 1714281807
transform 1 0 1204 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_646
timestamp 1714281807
transform 1 0 1204 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_647
timestamp 1714281807
transform 1 0 1132 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_648
timestamp 1714281807
transform 1 0 684 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_649
timestamp 1714281807
transform 1 0 684 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_650
timestamp 1714281807
transform 1 0 684 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_651
timestamp 1714281807
transform 1 0 2852 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_652
timestamp 1714281807
transform 1 0 2852 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_653
timestamp 1714281807
transform 1 0 2820 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_654
timestamp 1714281807
transform 1 0 2788 0 1 1785
box -2 -2 2 2
use M2_M1  M2_M1_655
timestamp 1714281807
transform 1 0 2788 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_656
timestamp 1714281807
transform 1 0 2788 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_657
timestamp 1714281807
transform 1 0 2788 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_658
timestamp 1714281807
transform 1 0 2732 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_659
timestamp 1714281807
transform 1 0 2724 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_660
timestamp 1714281807
transform 1 0 2716 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_661
timestamp 1714281807
transform 1 0 2572 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_662
timestamp 1714281807
transform 1 0 2556 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_663
timestamp 1714281807
transform 1 0 2516 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_664
timestamp 1714281807
transform 1 0 2396 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_665
timestamp 1714281807
transform 1 0 2220 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_666
timestamp 1714281807
transform 1 0 2204 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_667
timestamp 1714281807
transform 1 0 2108 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_668
timestamp 1714281807
transform 1 0 2108 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_669
timestamp 1714281807
transform 1 0 2092 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_670
timestamp 1714281807
transform 1 0 2068 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_671
timestamp 1714281807
transform 1 0 2020 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_672
timestamp 1714281807
transform 1 0 1996 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_673
timestamp 1714281807
transform 1 0 1996 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_674
timestamp 1714281807
transform 1 0 1988 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_675
timestamp 1714281807
transform 1 0 1956 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_676
timestamp 1714281807
transform 1 0 1956 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_677
timestamp 1714281807
transform 1 0 1844 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_678
timestamp 1714281807
transform 1 0 1708 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_679
timestamp 1714281807
transform 1 0 1676 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_680
timestamp 1714281807
transform 1 0 1596 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_681
timestamp 1714281807
transform 1 0 1564 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_682
timestamp 1714281807
transform 1 0 1516 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_683
timestamp 1714281807
transform 1 0 1500 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_684
timestamp 1714281807
transform 1 0 1348 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_685
timestamp 1714281807
transform 1 0 1236 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_686
timestamp 1714281807
transform 1 0 1188 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_687
timestamp 1714281807
transform 1 0 2860 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_688
timestamp 1714281807
transform 1 0 2852 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_689
timestamp 1714281807
transform 1 0 2836 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_690
timestamp 1714281807
transform 1 0 2820 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_691
timestamp 1714281807
transform 1 0 2812 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_692
timestamp 1714281807
transform 1 0 2812 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_693
timestamp 1714281807
transform 1 0 2772 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_694
timestamp 1714281807
transform 1 0 2724 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_695
timestamp 1714281807
transform 1 0 2684 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_696
timestamp 1714281807
transform 1 0 2636 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_697
timestamp 1714281807
transform 1 0 2620 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_698
timestamp 1714281807
transform 1 0 2580 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_699
timestamp 1714281807
transform 1 0 2508 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_700
timestamp 1714281807
transform 1 0 2500 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_701
timestamp 1714281807
transform 1 0 2492 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_702
timestamp 1714281807
transform 1 0 2468 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_703
timestamp 1714281807
transform 1 0 2420 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_704
timestamp 1714281807
transform 1 0 2396 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_705
timestamp 1714281807
transform 1 0 2388 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_706
timestamp 1714281807
transform 1 0 2284 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_707
timestamp 1714281807
transform 1 0 2268 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_708
timestamp 1714281807
transform 1 0 2252 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_709
timestamp 1714281807
transform 1 0 2236 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_710
timestamp 1714281807
transform 1 0 2092 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_711
timestamp 1714281807
transform 1 0 2076 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_712
timestamp 1714281807
transform 1 0 2052 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_713
timestamp 1714281807
transform 1 0 2020 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_714
timestamp 1714281807
transform 1 0 1612 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_715
timestamp 1714281807
transform 1 0 1604 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_716
timestamp 1714281807
transform 1 0 1564 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_717
timestamp 1714281807
transform 1 0 1548 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_718
timestamp 1714281807
transform 1 0 1524 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_719
timestamp 1714281807
transform 1 0 1468 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_720
timestamp 1714281807
transform 1 0 1468 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_721
timestamp 1714281807
transform 1 0 1452 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_722
timestamp 1714281807
transform 1 0 1060 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_723
timestamp 1714281807
transform 1 0 2684 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_724
timestamp 1714281807
transform 1 0 2628 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_725
timestamp 1714281807
transform 1 0 2572 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_726
timestamp 1714281807
transform 1 0 2556 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_727
timestamp 1714281807
transform 1 0 2460 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_728
timestamp 1714281807
transform 1 0 2420 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_729
timestamp 1714281807
transform 1 0 2412 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_730
timestamp 1714281807
transform 1 0 2404 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_731
timestamp 1714281807
transform 1 0 2228 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_732
timestamp 1714281807
transform 1 0 2076 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_733
timestamp 1714281807
transform 1 0 1964 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_734
timestamp 1714281807
transform 1 0 1804 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_735
timestamp 1714281807
transform 1 0 1788 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_736
timestamp 1714281807
transform 1 0 1308 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_737
timestamp 1714281807
transform 1 0 1068 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_738
timestamp 1714281807
transform 1 0 1068 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_739
timestamp 1714281807
transform 1 0 1036 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_740
timestamp 1714281807
transform 1 0 996 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_741
timestamp 1714281807
transform 1 0 1068 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_742
timestamp 1714281807
transform 1 0 1060 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_743
timestamp 1714281807
transform 1 0 1020 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_744
timestamp 1714281807
transform 1 0 1372 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_745
timestamp 1714281807
transform 1 0 1268 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_746
timestamp 1714281807
transform 1 0 1252 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_747
timestamp 1714281807
transform 1 0 1244 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_748
timestamp 1714281807
transform 1 0 1348 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_749
timestamp 1714281807
transform 1 0 1324 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_750
timestamp 1714281807
transform 1 0 1300 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_751
timestamp 1714281807
transform 1 0 1228 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_752
timestamp 1714281807
transform 1 0 1188 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_753
timestamp 1714281807
transform 1 0 2684 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_754
timestamp 1714281807
transform 1 0 2612 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_755
timestamp 1714281807
transform 1 0 2540 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_756
timestamp 1714281807
transform 1 0 2532 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_757
timestamp 1714281807
transform 1 0 2316 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_758
timestamp 1714281807
transform 1 0 2228 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_759
timestamp 1714281807
transform 1 0 2220 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_760
timestamp 1714281807
transform 1 0 2172 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_761
timestamp 1714281807
transform 1 0 1924 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_762
timestamp 1714281807
transform 1 0 1748 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_763
timestamp 1714281807
transform 1 0 1676 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_764
timestamp 1714281807
transform 1 0 1636 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_765
timestamp 1714281807
transform 1 0 1444 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_766
timestamp 1714281807
transform 1 0 1356 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_767
timestamp 1714281807
transform 1 0 1332 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_768
timestamp 1714281807
transform 1 0 1332 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_769
timestamp 1714281807
transform 1 0 1252 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_770
timestamp 1714281807
transform 1 0 1212 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_771
timestamp 1714281807
transform 1 0 1212 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_772
timestamp 1714281807
transform 1 0 1212 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_773
timestamp 1714281807
transform 1 0 1212 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_774
timestamp 1714281807
transform 1 0 1204 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_775
timestamp 1714281807
transform 1 0 1188 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_776
timestamp 1714281807
transform 1 0 1148 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_777
timestamp 1714281807
transform 1 0 1132 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_778
timestamp 1714281807
transform 1 0 1132 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_779
timestamp 1714281807
transform 1 0 812 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_780
timestamp 1714281807
transform 1 0 732 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_781
timestamp 1714281807
transform 1 0 556 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_782
timestamp 1714281807
transform 1 0 556 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_783
timestamp 1714281807
transform 1 0 412 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_784
timestamp 1714281807
transform 1 0 396 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_785
timestamp 1714281807
transform 1 0 372 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_786
timestamp 1714281807
transform 1 0 372 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_787
timestamp 1714281807
transform 1 0 1388 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_788
timestamp 1714281807
transform 1 0 1380 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_789
timestamp 1714281807
transform 1 0 1380 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_790
timestamp 1714281807
transform 1 0 1300 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_791
timestamp 1714281807
transform 1 0 1300 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_792
timestamp 1714281807
transform 1 0 1300 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_793
timestamp 1714281807
transform 1 0 1172 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_794
timestamp 1714281807
transform 1 0 1172 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_795
timestamp 1714281807
transform 1 0 1124 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_796
timestamp 1714281807
transform 1 0 1116 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_797
timestamp 1714281807
transform 1 0 1076 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_798
timestamp 1714281807
transform 1 0 1044 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_799
timestamp 1714281807
transform 1 0 1036 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_800
timestamp 1714281807
transform 1 0 2836 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_801
timestamp 1714281807
transform 1 0 2820 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_802
timestamp 1714281807
transform 1 0 2780 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_803
timestamp 1714281807
transform 1 0 2772 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_804
timestamp 1714281807
transform 1 0 2492 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_805
timestamp 1714281807
transform 1 0 2404 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_806
timestamp 1714281807
transform 1 0 2348 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_807
timestamp 1714281807
transform 1 0 2324 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_808
timestamp 1714281807
transform 1 0 2316 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_809
timestamp 1714281807
transform 1 0 2028 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_810
timestamp 1714281807
transform 1 0 1948 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_811
timestamp 1714281807
transform 1 0 1860 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_812
timestamp 1714281807
transform 1 0 1684 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_813
timestamp 1714281807
transform 1 0 1564 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_814
timestamp 1714281807
transform 1 0 1420 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_815
timestamp 1714281807
transform 1 0 1228 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_816
timestamp 1714281807
transform 1 0 1196 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_817
timestamp 1714281807
transform 1 0 1084 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_818
timestamp 1714281807
transform 1 0 2756 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_819
timestamp 1714281807
transform 1 0 2756 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_820
timestamp 1714281807
transform 1 0 2580 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_821
timestamp 1714281807
transform 1 0 2540 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_822
timestamp 1714281807
transform 1 0 2356 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_823
timestamp 1714281807
transform 1 0 2300 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_824
timestamp 1714281807
transform 1 0 2228 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_825
timestamp 1714281807
transform 1 0 2132 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_826
timestamp 1714281807
transform 1 0 1908 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_827
timestamp 1714281807
transform 1 0 1804 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_828
timestamp 1714281807
transform 1 0 1804 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_829
timestamp 1714281807
transform 1 0 1772 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_830
timestamp 1714281807
transform 1 0 1748 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_831
timestamp 1714281807
transform 1 0 1508 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_832
timestamp 1714281807
transform 1 0 1444 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_833
timestamp 1714281807
transform 1 0 1332 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_834
timestamp 1714281807
transform 1 0 1260 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_835
timestamp 1714281807
transform 1 0 1260 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_836
timestamp 1714281807
transform 1 0 2836 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_837
timestamp 1714281807
transform 1 0 2780 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_838
timestamp 1714281807
transform 1 0 2772 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_839
timestamp 1714281807
transform 1 0 2732 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_840
timestamp 1714281807
transform 1 0 2588 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_841
timestamp 1714281807
transform 1 0 2316 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_842
timestamp 1714281807
transform 1 0 2316 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_843
timestamp 1714281807
transform 1 0 2308 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_844
timestamp 1714281807
transform 1 0 2276 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_845
timestamp 1714281807
transform 1 0 2116 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_846
timestamp 1714281807
transform 1 0 1828 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_847
timestamp 1714281807
transform 1 0 1740 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_848
timestamp 1714281807
transform 1 0 1724 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_849
timestamp 1714281807
transform 1 0 1716 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_850
timestamp 1714281807
transform 1 0 1452 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_851
timestamp 1714281807
transform 1 0 1268 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_852
timestamp 1714281807
transform 1 0 1220 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_853
timestamp 1714281807
transform 1 0 1164 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_854
timestamp 1714281807
transform 1 0 1180 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_855
timestamp 1714281807
transform 1 0 980 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_856
timestamp 1714281807
transform 1 0 972 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_857
timestamp 1714281807
transform 1 0 884 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_858
timestamp 1714281807
transform 1 0 796 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_859
timestamp 1714281807
transform 1 0 572 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_860
timestamp 1714281807
transform 1 0 508 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_861
timestamp 1714281807
transform 1 0 460 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_862
timestamp 1714281807
transform 1 0 444 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_863
timestamp 1714281807
transform 1 0 404 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_864
timestamp 1714281807
transform 1 0 340 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_865
timestamp 1714281807
transform 1 0 316 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_866
timestamp 1714281807
transform 1 0 844 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_867
timestamp 1714281807
transform 1 0 788 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_868
timestamp 1714281807
transform 1 0 684 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_869
timestamp 1714281807
transform 1 0 620 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_870
timestamp 1714281807
transform 1 0 620 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_871
timestamp 1714281807
transform 1 0 564 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_872
timestamp 1714281807
transform 1 0 548 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_873
timestamp 1714281807
transform 1 0 476 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_874
timestamp 1714281807
transform 1 0 468 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_875
timestamp 1714281807
transform 1 0 412 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_876
timestamp 1714281807
transform 1 0 1020 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_877
timestamp 1714281807
transform 1 0 892 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_878
timestamp 1714281807
transform 1 0 1212 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_879
timestamp 1714281807
transform 1 0 972 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_880
timestamp 1714281807
transform 1 0 1132 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_881
timestamp 1714281807
transform 1 0 988 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_882
timestamp 1714281807
transform 1 0 1108 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_883
timestamp 1714281807
transform 1 0 1108 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_884
timestamp 1714281807
transform 1 0 1076 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_885
timestamp 1714281807
transform 1 0 948 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_886
timestamp 1714281807
transform 1 0 828 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_887
timestamp 1714281807
transform 1 0 756 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_888
timestamp 1714281807
transform 1 0 732 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_889
timestamp 1714281807
transform 1 0 548 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_890
timestamp 1714281807
transform 1 0 492 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_891
timestamp 1714281807
transform 1 0 492 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_892
timestamp 1714281807
transform 1 0 428 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_893
timestamp 1714281807
transform 1 0 260 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_894
timestamp 1714281807
transform 1 0 260 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_895
timestamp 1714281807
transform 1 0 1052 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_896
timestamp 1714281807
transform 1 0 1012 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_897
timestamp 1714281807
transform 1 0 900 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_898
timestamp 1714281807
transform 1 0 1332 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_899
timestamp 1714281807
transform 1 0 1292 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_900
timestamp 1714281807
transform 1 0 1324 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_901
timestamp 1714281807
transform 1 0 1188 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_902
timestamp 1714281807
transform 1 0 1236 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_903
timestamp 1714281807
transform 1 0 1036 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_904
timestamp 1714281807
transform 1 0 1212 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_905
timestamp 1714281807
transform 1 0 1012 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_906
timestamp 1714281807
transform 1 0 548 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_907
timestamp 1714281807
transform 1 0 548 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_908
timestamp 1714281807
transform 1 0 516 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_909
timestamp 1714281807
transform 1 0 396 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_910
timestamp 1714281807
transform 1 0 628 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_911
timestamp 1714281807
transform 1 0 380 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_912
timestamp 1714281807
transform 1 0 644 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_913
timestamp 1714281807
transform 1 0 500 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_914
timestamp 1714281807
transform 1 0 996 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_915
timestamp 1714281807
transform 1 0 916 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_916
timestamp 1714281807
transform 1 0 860 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_917
timestamp 1714281807
transform 1 0 852 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_918
timestamp 1714281807
transform 1 0 1100 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_919
timestamp 1714281807
transform 1 0 956 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_920
timestamp 1714281807
transform 1 0 1148 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_921
timestamp 1714281807
transform 1 0 1100 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_922
timestamp 1714281807
transform 1 0 972 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_923
timestamp 1714281807
transform 1 0 924 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_924
timestamp 1714281807
transform 1 0 860 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_925
timestamp 1714281807
transform 1 0 1028 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_926
timestamp 1714281807
transform 1 0 988 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_927
timestamp 1714281807
transform 1 0 956 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_928
timestamp 1714281807
transform 1 0 1196 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_929
timestamp 1714281807
transform 1 0 1148 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_930
timestamp 1714281807
transform 1 0 1116 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_931
timestamp 1714281807
transform 1 0 1244 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_932
timestamp 1714281807
transform 1 0 1188 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_933
timestamp 1714281807
transform 1 0 1156 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_934
timestamp 1714281807
transform 1 0 484 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_935
timestamp 1714281807
transform 1 0 484 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_936
timestamp 1714281807
transform 1 0 372 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_937
timestamp 1714281807
transform 1 0 356 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_938
timestamp 1714281807
transform 1 0 300 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_939
timestamp 1714281807
transform 1 0 268 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_940
timestamp 1714281807
transform 1 0 372 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_941
timestamp 1714281807
transform 1 0 316 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_942
timestamp 1714281807
transform 1 0 284 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_943
timestamp 1714281807
transform 1 0 516 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_944
timestamp 1714281807
transform 1 0 516 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_945
timestamp 1714281807
transform 1 0 476 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_946
timestamp 1714281807
transform 1 0 436 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_947
timestamp 1714281807
transform 1 0 1084 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_948
timestamp 1714281807
transform 1 0 1084 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_949
timestamp 1714281807
transform 1 0 932 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_950
timestamp 1714281807
transform 1 0 796 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_951
timestamp 1714281807
transform 1 0 772 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_952
timestamp 1714281807
transform 1 0 796 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_953
timestamp 1714281807
transform 1 0 676 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_954
timestamp 1714281807
transform 1 0 596 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_955
timestamp 1714281807
transform 1 0 868 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_956
timestamp 1714281807
transform 1 0 700 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_957
timestamp 1714281807
transform 1 0 548 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_958
timestamp 1714281807
transform 1 0 1100 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_959
timestamp 1714281807
transform 1 0 892 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_960
timestamp 1714281807
transform 1 0 820 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_961
timestamp 1714281807
transform 1 0 788 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_962
timestamp 1714281807
transform 1 0 724 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_963
timestamp 1714281807
transform 1 0 660 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_964
timestamp 1714281807
transform 1 0 620 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_965
timestamp 1714281807
transform 1 0 572 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_966
timestamp 1714281807
transform 1 0 540 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_967
timestamp 1714281807
transform 1 0 564 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_968
timestamp 1714281807
transform 1 0 556 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_969
timestamp 1714281807
transform 1 0 380 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_970
timestamp 1714281807
transform 1 0 676 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_971
timestamp 1714281807
transform 1 0 532 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_972
timestamp 1714281807
transform 1 0 396 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_973
timestamp 1714281807
transform 1 0 308 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_974
timestamp 1714281807
transform 1 0 212 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_975
timestamp 1714281807
transform 1 0 284 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_976
timestamp 1714281807
transform 1 0 228 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_977
timestamp 1714281807
transform 1 0 228 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_978
timestamp 1714281807
transform 1 0 300 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_979
timestamp 1714281807
transform 1 0 276 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_980
timestamp 1714281807
transform 1 0 276 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_981
timestamp 1714281807
transform 1 0 460 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_982
timestamp 1714281807
transform 1 0 452 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_983
timestamp 1714281807
transform 1 0 452 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_984
timestamp 1714281807
transform 1 0 876 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_985
timestamp 1714281807
transform 1 0 644 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_986
timestamp 1714281807
transform 1 0 644 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_987
timestamp 1714281807
transform 1 0 972 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_988
timestamp 1714281807
transform 1 0 820 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_989
timestamp 1714281807
transform 1 0 1164 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_990
timestamp 1714281807
transform 1 0 1132 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_991
timestamp 1714281807
transform 1 0 1076 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_992
timestamp 1714281807
transform 1 0 1172 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_993
timestamp 1714281807
transform 1 0 1092 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_994
timestamp 1714281807
transform 1 0 1020 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_995
timestamp 1714281807
transform 1 0 956 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_996
timestamp 1714281807
transform 1 0 468 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_997
timestamp 1714281807
transform 1 0 420 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_998
timestamp 1714281807
transform 1 0 420 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_999
timestamp 1714281807
transform 1 0 396 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1000
timestamp 1714281807
transform 1 0 380 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_1001
timestamp 1714281807
transform 1 0 1140 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1002
timestamp 1714281807
transform 1 0 1108 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1003
timestamp 1714281807
transform 1 0 1100 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1004
timestamp 1714281807
transform 1 0 628 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1005
timestamp 1714281807
transform 1 0 580 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1006
timestamp 1714281807
transform 1 0 580 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1007
timestamp 1714281807
transform 1 0 540 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1008
timestamp 1714281807
transform 1 0 428 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_1009
timestamp 1714281807
transform 1 0 308 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1010
timestamp 1714281807
transform 1 0 244 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1011
timestamp 1714281807
transform 1 0 1036 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1012
timestamp 1714281807
transform 1 0 932 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1013
timestamp 1714281807
transform 1 0 812 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1014
timestamp 1714281807
transform 1 0 812 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1015
timestamp 1714281807
transform 1 0 684 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_1016
timestamp 1714281807
transform 1 0 660 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1017
timestamp 1714281807
transform 1 0 652 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1018
timestamp 1714281807
transform 1 0 532 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1019
timestamp 1714281807
transform 1 0 444 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1020
timestamp 1714281807
transform 1 0 420 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1021
timestamp 1714281807
transform 1 0 372 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1022
timestamp 1714281807
transform 1 0 260 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1023
timestamp 1714281807
transform 1 0 212 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1024
timestamp 1714281807
transform 1 0 204 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1025
timestamp 1714281807
transform 1 0 836 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_1026
timestamp 1714281807
transform 1 0 812 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1027
timestamp 1714281807
transform 1 0 676 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_1028
timestamp 1714281807
transform 1 0 652 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1029
timestamp 1714281807
transform 1 0 436 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1030
timestamp 1714281807
transform 1 0 316 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_1031
timestamp 1714281807
transform 1 0 524 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1032
timestamp 1714281807
transform 1 0 492 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_1033
timestamp 1714281807
transform 1 0 724 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1034
timestamp 1714281807
transform 1 0 692 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_1035
timestamp 1714281807
transform 1 0 884 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1036
timestamp 1714281807
transform 1 0 860 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_1037
timestamp 1714281807
transform 1 0 980 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1038
timestamp 1714281807
transform 1 0 948 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1039
timestamp 1714281807
transform 1 0 932 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1040
timestamp 1714281807
transform 1 0 868 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1041
timestamp 1714281807
transform 1 0 916 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1042
timestamp 1714281807
transform 1 0 764 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1043
timestamp 1714281807
transform 1 0 868 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1044
timestamp 1714281807
transform 1 0 868 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1045
timestamp 1714281807
transform 1 0 1044 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1046
timestamp 1714281807
transform 1 0 964 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1047
timestamp 1714281807
transform 1 0 1196 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1048
timestamp 1714281807
transform 1 0 1124 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1049
timestamp 1714281807
transform 1 0 1252 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1050
timestamp 1714281807
transform 1 0 1164 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1051
timestamp 1714281807
transform 1 0 1092 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1052
timestamp 1714281807
transform 1 0 996 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1053
timestamp 1714281807
transform 1 0 780 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1054
timestamp 1714281807
transform 1 0 748 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1055
timestamp 1714281807
transform 1 0 612 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1056
timestamp 1714281807
transform 1 0 612 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1057
timestamp 1714281807
transform 1 0 628 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1058
timestamp 1714281807
transform 1 0 556 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1059
timestamp 1714281807
transform 1 0 876 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1060
timestamp 1714281807
transform 1 0 836 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1061
timestamp 1714281807
transform 1 0 716 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1062
timestamp 1714281807
transform 1 0 676 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1063
timestamp 1714281807
transform 1 0 548 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1064
timestamp 1714281807
transform 1 0 492 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1065
timestamp 1714281807
transform 1 0 388 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1066
timestamp 1714281807
transform 1 0 284 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1067
timestamp 1714281807
transform 1 0 524 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1068
timestamp 1714281807
transform 1 0 396 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1069
timestamp 1714281807
transform 1 0 276 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1070
timestamp 1714281807
transform 1 0 236 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1071
timestamp 1714281807
transform 1 0 292 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1072
timestamp 1714281807
transform 1 0 212 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1073
timestamp 1714281807
transform 1 0 444 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1074
timestamp 1714281807
transform 1 0 380 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1075
timestamp 1714281807
transform 1 0 220 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1076
timestamp 1714281807
transform 1 0 220 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1077
timestamp 1714281807
transform 1 0 268 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1078
timestamp 1714281807
transform 1 0 156 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1079
timestamp 1714281807
transform 1 0 292 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1080
timestamp 1714281807
transform 1 0 180 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1081
timestamp 1714281807
transform 1 0 468 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1082
timestamp 1714281807
transform 1 0 380 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1083
timestamp 1714281807
transform 1 0 676 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1084
timestamp 1714281807
transform 1 0 604 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1085
timestamp 1714281807
transform 1 0 836 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1086
timestamp 1714281807
transform 1 0 804 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1087
timestamp 1714281807
transform 1 0 1092 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1088
timestamp 1714281807
transform 1 0 1084 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1089
timestamp 1714281807
transform 1 0 996 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1090
timestamp 1714281807
transform 1 0 964 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1091
timestamp 1714281807
transform 1 0 1412 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1092
timestamp 1714281807
transform 1 0 1276 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1093
timestamp 1714281807
transform 1 0 2204 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1094
timestamp 1714281807
transform 1 0 2140 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1095
timestamp 1714281807
transform 1 0 2204 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1096
timestamp 1714281807
transform 1 0 2164 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1097
timestamp 1714281807
transform 1 0 1892 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1098
timestamp 1714281807
transform 1 0 1892 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1099
timestamp 1714281807
transform 1 0 2068 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1100
timestamp 1714281807
transform 1 0 2020 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1101
timestamp 1714281807
transform 1 0 2116 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1102
timestamp 1714281807
transform 1 0 2076 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1103
timestamp 1714281807
transform 1 0 2116 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1104
timestamp 1714281807
transform 1 0 2116 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1105
timestamp 1714281807
transform 1 0 1556 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1106
timestamp 1714281807
transform 1 0 1516 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1107
timestamp 1714281807
transform 1 0 1500 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1108
timestamp 1714281807
transform 1 0 1460 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1109
timestamp 1714281807
transform 1 0 1564 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1110
timestamp 1714281807
transform 1 0 1564 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_1111
timestamp 1714281807
transform 1 0 1556 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1112
timestamp 1714281807
transform 1 0 1516 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1113
timestamp 1714281807
transform 1 0 1692 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1114
timestamp 1714281807
transform 1 0 1652 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1115
timestamp 1714281807
transform 1 0 1548 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1116
timestamp 1714281807
transform 1 0 1508 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1117
timestamp 1714281807
transform 1 0 1660 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1118
timestamp 1714281807
transform 1 0 1612 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1119
timestamp 1714281807
transform 1 0 2108 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1120
timestamp 1714281807
transform 1 0 2068 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1121
timestamp 1714281807
transform 1 0 2044 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1122
timestamp 1714281807
transform 1 0 2004 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1123
timestamp 1714281807
transform 1 0 2228 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1124
timestamp 1714281807
transform 1 0 2156 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1125
timestamp 1714281807
transform 1 0 2196 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1126
timestamp 1714281807
transform 1 0 2196 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_1127
timestamp 1714281807
transform 1 0 1868 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1128
timestamp 1714281807
transform 1 0 1868 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1129
timestamp 1714281807
transform 1 0 2612 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1130
timestamp 1714281807
transform 1 0 2604 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_1131
timestamp 1714281807
transform 1 0 2604 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1132
timestamp 1714281807
transform 1 0 2564 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1133
timestamp 1714281807
transform 1 0 2380 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1134
timestamp 1714281807
transform 1 0 2332 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1135
timestamp 1714281807
transform 1 0 2884 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1136
timestamp 1714281807
transform 1 0 2844 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1137
timestamp 1714281807
transform 1 0 2892 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1138
timestamp 1714281807
transform 1 0 2852 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1139
timestamp 1714281807
transform 1 0 2812 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1140
timestamp 1714281807
transform 1 0 2772 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1141
timestamp 1714281807
transform 1 0 2380 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1142
timestamp 1714281807
transform 1 0 2340 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1143
timestamp 1714281807
transform 1 0 2572 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1144
timestamp 1714281807
transform 1 0 2532 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1145
timestamp 1714281807
transform 1 0 2228 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1146
timestamp 1714281807
transform 1 0 2172 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1147
timestamp 1714281807
transform 1 0 2812 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1148
timestamp 1714281807
transform 1 0 2772 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1149
timestamp 1714281807
transform 1 0 2908 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1150
timestamp 1714281807
transform 1 0 2868 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1151
timestamp 1714281807
transform 1 0 2564 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1152
timestamp 1714281807
transform 1 0 2524 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1153
timestamp 1714281807
transform 1 0 1644 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1154
timestamp 1714281807
transform 1 0 1604 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1155
timestamp 1714281807
transform 1 0 1684 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1156
timestamp 1714281807
transform 1 0 1636 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1157
timestamp 1714281807
transform 1 0 1652 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1158
timestamp 1714281807
transform 1 0 1612 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1159
timestamp 1714281807
transform 1 0 2908 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1160
timestamp 1714281807
transform 1 0 2868 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1161
timestamp 1714281807
transform 1 0 2852 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1162
timestamp 1714281807
transform 1 0 2796 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1163
timestamp 1714281807
transform 1 0 2500 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_1164
timestamp 1714281807
transform 1 0 2500 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1165
timestamp 1714281807
transform 1 0 2020 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1166
timestamp 1714281807
transform 1 0 2020 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1167
timestamp 1714281807
transform 1 0 2028 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1168
timestamp 1714281807
transform 1 0 1988 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1169
timestamp 1714281807
transform 1 0 1788 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1170
timestamp 1714281807
transform 1 0 1772 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1171
timestamp 1714281807
transform 1 0 2380 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_1172
timestamp 1714281807
transform 1 0 2380 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1173
timestamp 1714281807
transform 1 0 2276 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1174
timestamp 1714281807
transform 1 0 2276 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1175
timestamp 1714281807
transform 1 0 2124 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1176
timestamp 1714281807
transform 1 0 2124 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1177
timestamp 1714281807
transform 1 0 2908 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1178
timestamp 1714281807
transform 1 0 2868 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1179
timestamp 1714281807
transform 1 0 2900 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1180
timestamp 1714281807
transform 1 0 2860 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1181
timestamp 1714281807
transform 1 0 2900 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1182
timestamp 1714281807
transform 1 0 2860 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1183
timestamp 1714281807
transform 1 0 2244 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1184
timestamp 1714281807
transform 1 0 2204 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1185
timestamp 1714281807
transform 1 0 2044 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1186
timestamp 1714281807
transform 1 0 2044 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1187
timestamp 1714281807
transform 1 0 2164 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1188
timestamp 1714281807
transform 1 0 2116 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1189
timestamp 1714281807
transform 1 0 1644 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1190
timestamp 1714281807
transform 1 0 1604 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1191
timestamp 1714281807
transform 1 0 1612 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1192
timestamp 1714281807
transform 1 0 1564 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1193
timestamp 1714281807
transform 1 0 1748 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1194
timestamp 1714281807
transform 1 0 1748 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1195
timestamp 1714281807
transform 1 0 1780 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1196
timestamp 1714281807
transform 1 0 1780 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1197
timestamp 1714281807
transform 1 0 1684 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1198
timestamp 1714281807
transform 1 0 1684 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1199
timestamp 1714281807
transform 1 0 1796 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1200
timestamp 1714281807
transform 1 0 1796 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1201
timestamp 1714281807
transform 1 0 1012 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1202
timestamp 1714281807
transform 1 0 972 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1203
timestamp 1714281807
transform 1 0 1060 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1204
timestamp 1714281807
transform 1 0 964 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1205
timestamp 1714281807
transform 1 0 1100 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1206
timestamp 1714281807
transform 1 0 1100 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1207
timestamp 1714281807
transform 1 0 1012 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1208
timestamp 1714281807
transform 1 0 972 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1209
timestamp 1714281807
transform 1 0 980 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_1210
timestamp 1714281807
transform 1 0 980 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1211
timestamp 1714281807
transform 1 0 1156 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1212
timestamp 1714281807
transform 1 0 1108 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1213
timestamp 1714281807
transform 1 0 1516 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1214
timestamp 1714281807
transform 1 0 1476 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1215
timestamp 1714281807
transform 1 0 1676 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1216
timestamp 1714281807
transform 1 0 1636 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1217
timestamp 1714281807
transform 1 0 1340 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1218
timestamp 1714281807
transform 1 0 1300 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1219
timestamp 1714281807
transform 1 0 2156 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1220
timestamp 1714281807
transform 1 0 2116 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1221
timestamp 1714281807
transform 1 0 1988 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1222
timestamp 1714281807
transform 1 0 1948 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1223
timestamp 1714281807
transform 1 0 1844 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1224
timestamp 1714281807
transform 1 0 1796 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1225
timestamp 1714281807
transform 1 0 2508 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1226
timestamp 1714281807
transform 1 0 2468 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1227
timestamp 1714281807
transform 1 0 2652 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1228
timestamp 1714281807
transform 1 0 2612 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1229
timestamp 1714281807
transform 1 0 2332 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1230
timestamp 1714281807
transform 1 0 2292 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1231
timestamp 1714281807
transform 1 0 2940 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1232
timestamp 1714281807
transform 1 0 2900 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1233
timestamp 1714281807
transform 1 0 2940 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1234
timestamp 1714281807
transform 1 0 2900 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1235
timestamp 1714281807
transform 1 0 2788 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1236
timestamp 1714281807
transform 1 0 2748 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1237
timestamp 1714281807
transform 1 0 2524 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1238
timestamp 1714281807
transform 1 0 2524 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1239
timestamp 1714281807
transform 1 0 2508 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1240
timestamp 1714281807
transform 1 0 2468 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1241
timestamp 1714281807
transform 1 0 2652 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1242
timestamp 1714281807
transform 1 0 2612 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1243
timestamp 1714281807
transform 1 0 2884 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1244
timestamp 1714281807
transform 1 0 2884 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1245
timestamp 1714281807
transform 1 0 2820 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1246
timestamp 1714281807
transform 1 0 2780 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1247
timestamp 1714281807
transform 1 0 2692 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1248
timestamp 1714281807
transform 1 0 2644 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1249
timestamp 1714281807
transform 1 0 1636 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1250
timestamp 1714281807
transform 1 0 1596 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1251
timestamp 1714281807
transform 1 0 1684 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1252
timestamp 1714281807
transform 1 0 1644 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1253
timestamp 1714281807
transform 1 0 1604 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1254
timestamp 1714281807
transform 1 0 1564 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1255
timestamp 1714281807
transform 1 0 2860 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1256
timestamp 1714281807
transform 1 0 2836 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1257
timestamp 1714281807
transform 1 0 2716 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1258
timestamp 1714281807
transform 1 0 2716 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1259
timestamp 1714281807
transform 1 0 2612 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1260
timestamp 1714281807
transform 1 0 2612 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1261
timestamp 1714281807
transform 1 0 2052 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1262
timestamp 1714281807
transform 1 0 2020 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1263
timestamp 1714281807
transform 1 0 1916 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1264
timestamp 1714281807
transform 1 0 1876 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1265
timestamp 1714281807
transform 1 0 1772 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1266
timestamp 1714281807
transform 1 0 1724 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1267
timestamp 1714281807
transform 1 0 2500 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1268
timestamp 1714281807
transform 1 0 2444 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1269
timestamp 1714281807
transform 1 0 2332 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1270
timestamp 1714281807
transform 1 0 2292 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1271
timestamp 1714281807
transform 1 0 2172 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1272
timestamp 1714281807
transform 1 0 2124 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1273
timestamp 1714281807
transform 1 0 2612 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1274
timestamp 1714281807
transform 1 0 2572 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1275
timestamp 1714281807
transform 1 0 2572 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1276
timestamp 1714281807
transform 1 0 2532 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1277
timestamp 1714281807
transform 1 0 2668 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1278
timestamp 1714281807
transform 1 0 2628 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1279
timestamp 1714281807
transform 1 0 2532 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1280
timestamp 1714281807
transform 1 0 2492 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1281
timestamp 1714281807
transform 1 0 2556 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1282
timestamp 1714281807
transform 1 0 2540 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1283
timestamp 1714281807
transform 1 0 2516 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1284
timestamp 1714281807
transform 1 0 2428 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1285
timestamp 1714281807
transform 1 0 2828 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1286
timestamp 1714281807
transform 1 0 2812 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1287
timestamp 1714281807
transform 1 0 2732 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1288
timestamp 1714281807
transform 1 0 2708 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1289
timestamp 1714281807
transform 1 0 2836 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1290
timestamp 1714281807
transform 1 0 2820 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1291
timestamp 1714281807
transform 1 0 2748 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1292
timestamp 1714281807
transform 1 0 2724 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1293
timestamp 1714281807
transform 1 0 2844 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1294
timestamp 1714281807
transform 1 0 2828 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1295
timestamp 1714281807
transform 1 0 2764 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1296
timestamp 1714281807
transform 1 0 2732 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1297
timestamp 1714281807
transform 1 0 1420 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1298
timestamp 1714281807
transform 1 0 1420 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1299
timestamp 1714281807
transform 1 0 1420 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1300
timestamp 1714281807
transform 1 0 1380 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1301
timestamp 1714281807
transform 1 0 1044 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1302
timestamp 1714281807
transform 1 0 1044 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1303
timestamp 1714281807
transform 1 0 1492 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1304
timestamp 1714281807
transform 1 0 1452 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1305
timestamp 1714281807
transform 1 0 1420 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1306
timestamp 1714281807
transform 1 0 1372 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1307
timestamp 1714281807
transform 1 0 836 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1308
timestamp 1714281807
transform 1 0 796 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1309
timestamp 1714281807
transform 1 0 748 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1310
timestamp 1714281807
transform 1 0 732 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1311
timestamp 1714281807
transform 1 0 1452 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1312
timestamp 1714281807
transform 1 0 1452 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1313
timestamp 1714281807
transform 1 0 956 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1314
timestamp 1714281807
transform 1 0 956 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1315
timestamp 1714281807
transform 1 0 804 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1316
timestamp 1714281807
transform 1 0 764 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1317
timestamp 1714281807
transform 1 0 188 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1318
timestamp 1714281807
transform 1 0 148 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1319
timestamp 1714281807
transform 1 0 156 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1320
timestamp 1714281807
transform 1 0 156 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1321
timestamp 1714281807
transform 1 0 364 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1322
timestamp 1714281807
transform 1 0 356 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1323
timestamp 1714281807
transform 1 0 348 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1324
timestamp 1714281807
transform 1 0 268 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1325
timestamp 1714281807
transform 1 0 284 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1326
timestamp 1714281807
transform 1 0 284 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1327
timestamp 1714281807
transform 1 0 188 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1328
timestamp 1714281807
transform 1 0 188 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1329
timestamp 1714281807
transform 1 0 252 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1330
timestamp 1714281807
transform 1 0 252 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_1331
timestamp 1714281807
transform 1 0 364 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1332
timestamp 1714281807
transform 1 0 324 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1333
timestamp 1714281807
transform 1 0 540 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1334
timestamp 1714281807
transform 1 0 540 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1335
timestamp 1714281807
transform 1 0 292 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_1336
timestamp 1714281807
transform 1 0 292 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1337
timestamp 1714281807
transform 1 0 2220 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1338
timestamp 1714281807
transform 1 0 2116 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1339
timestamp 1714281807
transform 1 0 2116 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1340
timestamp 1714281807
transform 1 0 2124 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1341
timestamp 1714281807
transform 1 0 2100 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1342
timestamp 1714281807
transform 1 0 2740 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1343
timestamp 1714281807
transform 1 0 2724 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1344
timestamp 1714281807
transform 1 0 2676 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1345
timestamp 1714281807
transform 1 0 2652 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1346
timestamp 1714281807
transform 1 0 2860 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1347
timestamp 1714281807
transform 1 0 2836 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1348
timestamp 1714281807
transform 1 0 2748 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1349
timestamp 1714281807
transform 1 0 2812 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1350
timestamp 1714281807
transform 1 0 2796 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1351
timestamp 1714281807
transform 1 0 2748 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1352
timestamp 1714281807
transform 1 0 2740 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1353
timestamp 1714281807
transform 1 0 2132 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1354
timestamp 1714281807
transform 1 0 2116 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1355
timestamp 1714281807
transform 1 0 2284 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1356
timestamp 1714281807
transform 1 0 2284 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1357
timestamp 1714281807
transform 1 0 2204 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1358
timestamp 1714281807
transform 1 0 2412 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1359
timestamp 1714281807
transform 1 0 2412 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1360
timestamp 1714281807
transform 1 0 2332 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1361
timestamp 1714281807
transform 1 0 2748 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1362
timestamp 1714281807
transform 1 0 2708 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1363
timestamp 1714281807
transform 1 0 2708 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1364
timestamp 1714281807
transform 1 0 2652 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1365
timestamp 1714281807
transform 1 0 2644 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1366
timestamp 1714281807
transform 1 0 2884 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1367
timestamp 1714281807
transform 1 0 2884 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1368
timestamp 1714281807
transform 1 0 2852 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1369
timestamp 1714281807
transform 1 0 2836 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1370
timestamp 1714281807
transform 1 0 2828 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1371
timestamp 1714281807
transform 1 0 2868 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1372
timestamp 1714281807
transform 1 0 2860 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1373
timestamp 1714281807
transform 1 0 2780 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1374
timestamp 1714281807
transform 1 0 2660 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1375
timestamp 1714281807
transform 1 0 2596 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1376
timestamp 1714281807
transform 1 0 2380 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1377
timestamp 1714281807
transform 1 0 2228 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1378
timestamp 1714281807
transform 1 0 2140 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1379
timestamp 1714281807
transform 1 0 2436 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1380
timestamp 1714281807
transform 1 0 2436 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1381
timestamp 1714281807
transform 1 0 2420 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1382
timestamp 1714281807
transform 1 0 2332 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1383
timestamp 1714281807
transform 1 0 2524 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1384
timestamp 1714281807
transform 1 0 2364 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1385
timestamp 1714281807
transform 1 0 2364 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1386
timestamp 1714281807
transform 1 0 2324 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1387
timestamp 1714281807
transform 1 0 2316 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1388
timestamp 1714281807
transform 1 0 2700 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1389
timestamp 1714281807
transform 1 0 2692 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1390
timestamp 1714281807
transform 1 0 2660 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1391
timestamp 1714281807
transform 1 0 2628 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1392
timestamp 1714281807
transform 1 0 2852 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1393
timestamp 1714281807
transform 1 0 2852 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1394
timestamp 1714281807
transform 1 0 2828 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1395
timestamp 1714281807
transform 1 0 2796 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1396
timestamp 1714281807
transform 1 0 2796 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1397
timestamp 1714281807
transform 1 0 2900 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1398
timestamp 1714281807
transform 1 0 2884 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1399
timestamp 1714281807
transform 1 0 2852 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1400
timestamp 1714281807
transform 1 0 2836 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1401
timestamp 1714281807
transform 1 0 1540 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1402
timestamp 1714281807
transform 1 0 1524 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1403
timestamp 1714281807
transform 1 0 1492 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1404
timestamp 1714281807
transform 1 0 1484 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1405
timestamp 1714281807
transform 1 0 1444 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1406
timestamp 1714281807
transform 1 0 1636 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1407
timestamp 1714281807
transform 1 0 1572 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1408
timestamp 1714281807
transform 1 0 1372 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1409
timestamp 1714281807
transform 1 0 1300 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1410
timestamp 1714281807
transform 1 0 1580 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1411
timestamp 1714281807
transform 1 0 1508 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1412
timestamp 1714281807
transform 1 0 1356 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1413
timestamp 1714281807
transform 1 0 1756 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1414
timestamp 1714281807
transform 1 0 1732 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1415
timestamp 1714281807
transform 1 0 1972 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1416
timestamp 1714281807
transform 1 0 1876 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1417
timestamp 1714281807
transform 1 0 2036 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1418
timestamp 1714281807
transform 1 0 1972 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1419
timestamp 1714281807
transform 1 0 1956 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1420
timestamp 1714281807
transform 1 0 2636 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1421
timestamp 1714281807
transform 1 0 2620 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1422
timestamp 1714281807
transform 1 0 2596 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1423
timestamp 1714281807
transform 1 0 2572 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1424
timestamp 1714281807
transform 1 0 2532 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1425
timestamp 1714281807
transform 1 0 2508 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1426
timestamp 1714281807
transform 1 0 2708 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1427
timestamp 1714281807
transform 1 0 2692 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1428
timestamp 1714281807
transform 1 0 2636 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1429
timestamp 1714281807
transform 1 0 2892 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1430
timestamp 1714281807
transform 1 0 2876 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1431
timestamp 1714281807
transform 1 0 2836 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1432
timestamp 1714281807
transform 1 0 2828 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1433
timestamp 1714281807
transform 1 0 2804 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1434
timestamp 1714281807
transform 1 0 1804 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1435
timestamp 1714281807
transform 1 0 1804 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1436
timestamp 1714281807
transform 1 0 1804 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1437
timestamp 1714281807
transform 1 0 1764 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1438
timestamp 1714281807
transform 1 0 1916 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1439
timestamp 1714281807
transform 1 0 1860 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1440
timestamp 1714281807
transform 1 0 1860 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1441
timestamp 1714281807
transform 1 0 1860 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1442
timestamp 1714281807
transform 1 0 2076 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1443
timestamp 1714281807
transform 1 0 2028 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1444
timestamp 1714281807
transform 1 0 1956 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1445
timestamp 1714281807
transform 1 0 1948 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1446
timestamp 1714281807
transform 1 0 2108 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1447
timestamp 1714281807
transform 1 0 2100 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1448
timestamp 1714281807
transform 1 0 2100 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1449
timestamp 1714281807
transform 1 0 2060 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1450
timestamp 1714281807
transform 1 0 2284 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1451
timestamp 1714281807
transform 1 0 2284 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1452
timestamp 1714281807
transform 1 0 2220 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1453
timestamp 1714281807
transform 1 0 2220 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1454
timestamp 1714281807
transform 1 0 2436 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1455
timestamp 1714281807
transform 1 0 2404 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1456
timestamp 1714281807
transform 1 0 2348 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1457
timestamp 1714281807
transform 1 0 2348 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1458
timestamp 1714281807
transform 1 0 2708 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1459
timestamp 1714281807
transform 1 0 2700 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1460
timestamp 1714281807
transform 1 0 2676 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1461
timestamp 1714281807
transform 1 0 2868 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1462
timestamp 1714281807
transform 1 0 2844 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1463
timestamp 1714281807
transform 1 0 2804 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1464
timestamp 1714281807
transform 1 0 2628 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1465
timestamp 1714281807
transform 1 0 2844 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1466
timestamp 1714281807
transform 1 0 2844 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1467
timestamp 1714281807
transform 1 0 2788 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1468
timestamp 1714281807
transform 1 0 2652 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1469
timestamp 1714281807
transform 1 0 2636 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1470
timestamp 1714281807
transform 1 0 2524 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1471
timestamp 1714281807
transform 1 0 2516 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1472
timestamp 1714281807
transform 1 0 2492 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1473
timestamp 1714281807
transform 1 0 2836 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1474
timestamp 1714281807
transform 1 0 2820 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1475
timestamp 1714281807
transform 1 0 2780 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1476
timestamp 1714281807
transform 1 0 2644 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1477
timestamp 1714281807
transform 1 0 2732 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1478
timestamp 1714281807
transform 1 0 2716 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1479
timestamp 1714281807
transform 1 0 2636 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1480
timestamp 1714281807
transform 1 0 2612 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1481
timestamp 1714281807
transform 1 0 2540 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1482
timestamp 1714281807
transform 1 0 2540 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1483
timestamp 1714281807
transform 1 0 2468 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1484
timestamp 1714281807
transform 1 0 2788 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1485
timestamp 1714281807
transform 1 0 2620 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1486
timestamp 1714281807
transform 1 0 2596 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1487
timestamp 1714281807
transform 1 0 2828 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1488
timestamp 1714281807
transform 1 0 2804 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1489
timestamp 1714281807
transform 1 0 2692 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1490
timestamp 1714281807
transform 1 0 2436 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1491
timestamp 1714281807
transform 1 0 2420 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1492
timestamp 1714281807
transform 1 0 2332 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1493
timestamp 1714281807
transform 1 0 2588 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1494
timestamp 1714281807
transform 1 0 2548 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1495
timestamp 1714281807
transform 1 0 2372 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1496
timestamp 1714281807
transform 1 0 2308 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1497
timestamp 1714281807
transform 1 0 2476 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1498
timestamp 1714281807
transform 1 0 2348 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1499
timestamp 1714281807
transform 1 0 2332 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1500
timestamp 1714281807
transform 1 0 2276 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1501
timestamp 1714281807
transform 1 0 2244 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1502
timestamp 1714281807
transform 1 0 2132 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1503
timestamp 1714281807
transform 1 0 2116 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1504
timestamp 1714281807
transform 1 0 2084 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1505
timestamp 1714281807
transform 1 0 2084 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1506
timestamp 1714281807
transform 1 0 2116 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1507
timestamp 1714281807
transform 1 0 2108 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1508
timestamp 1714281807
transform 1 0 2092 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1509
timestamp 1714281807
transform 1 0 2124 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1510
timestamp 1714281807
transform 1 0 2028 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1511
timestamp 1714281807
transform 1 0 2004 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1512
timestamp 1714281807
transform 1 0 2052 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1513
timestamp 1714281807
transform 1 0 1964 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1514
timestamp 1714281807
transform 1 0 2012 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1515
timestamp 1714281807
transform 1 0 1988 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1516
timestamp 1714281807
transform 1 0 1564 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1517
timestamp 1714281807
transform 1 0 1532 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1518
timestamp 1714281807
transform 1 0 1444 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1519
timestamp 1714281807
transform 1 0 1452 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1520
timestamp 1714281807
transform 1 0 1380 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1521
timestamp 1714281807
transform 1 0 1492 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1522
timestamp 1714281807
transform 1 0 1476 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1523
timestamp 1714281807
transform 1 0 1444 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1524
timestamp 1714281807
transform 1 0 1444 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1525
timestamp 1714281807
transform 1 0 1588 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1526
timestamp 1714281807
transform 1 0 1572 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1527
timestamp 1714281807
transform 1 0 1524 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1528
timestamp 1714281807
transform 1 0 1500 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1529
timestamp 1714281807
transform 1 0 1644 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1530
timestamp 1714281807
transform 1 0 1628 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1531
timestamp 1714281807
transform 1 0 1572 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1532
timestamp 1714281807
transform 1 0 1548 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1533
timestamp 1714281807
transform 1 0 1580 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1534
timestamp 1714281807
transform 1 0 1492 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1535
timestamp 1714281807
transform 1 0 1420 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1536
timestamp 1714281807
transform 1 0 1484 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1537
timestamp 1714281807
transform 1 0 1396 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1538
timestamp 1714281807
transform 1 0 1652 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1539
timestamp 1714281807
transform 1 0 1652 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1540
timestamp 1714281807
transform 1 0 1492 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1541
timestamp 1714281807
transform 1 0 1396 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1542
timestamp 1714281807
transform 1 0 1972 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1543
timestamp 1714281807
transform 1 0 1956 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1544
timestamp 1714281807
transform 1 0 1900 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1545
timestamp 1714281807
transform 1 0 1860 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1546
timestamp 1714281807
transform 1 0 2052 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1547
timestamp 1714281807
transform 1 0 1964 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1548
timestamp 1714281807
transform 1 0 1724 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1549
timestamp 1714281807
transform 1 0 1724 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1550
timestamp 1714281807
transform 1 0 1860 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1551
timestamp 1714281807
transform 1 0 1780 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1552
timestamp 1714281807
transform 1 0 1780 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1553
timestamp 1714281807
transform 1 0 2220 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1554
timestamp 1714281807
transform 1 0 2172 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1555
timestamp 1714281807
transform 1 0 2092 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1556
timestamp 1714281807
transform 1 0 2124 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1557
timestamp 1714281807
transform 1 0 2020 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1558
timestamp 1714281807
transform 1 0 2020 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1559
timestamp 1714281807
transform 1 0 2324 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1560
timestamp 1714281807
transform 1 0 2316 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1561
timestamp 1714281807
transform 1 0 2548 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1562
timestamp 1714281807
transform 1 0 2540 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1563
timestamp 1714281807
transform 1 0 2476 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1564
timestamp 1714281807
transform 1 0 2572 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1565
timestamp 1714281807
transform 1 0 2508 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1566
timestamp 1714281807
transform 1 0 2404 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1567
timestamp 1714281807
transform 1 0 2260 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1568
timestamp 1714281807
transform 1 0 2260 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1569
timestamp 1714281807
transform 1 0 2500 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1570
timestamp 1714281807
transform 1 0 2468 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1571
timestamp 1714281807
transform 1 0 2444 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1572
timestamp 1714281807
transform 1 0 2428 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1573
timestamp 1714281807
transform 1 0 2420 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1574
timestamp 1714281807
transform 1 0 2380 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1575
timestamp 1714281807
transform 1 0 2380 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1576
timestamp 1714281807
transform 1 0 980 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1577
timestamp 1714281807
transform 1 0 972 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1578
timestamp 1714281807
transform 1 0 700 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1579
timestamp 1714281807
transform 1 0 532 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1580
timestamp 1714281807
transform 1 0 612 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1581
timestamp 1714281807
transform 1 0 516 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1582
timestamp 1714281807
transform 1 0 908 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1583
timestamp 1714281807
transform 1 0 764 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1584
timestamp 1714281807
transform 1 0 732 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1585
timestamp 1714281807
transform 1 0 676 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1586
timestamp 1714281807
transform 1 0 1004 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1587
timestamp 1714281807
transform 1 0 948 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1588
timestamp 1714281807
transform 1 0 932 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1589
timestamp 1714281807
transform 1 0 932 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1590
timestamp 1714281807
transform 1 0 604 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1591
timestamp 1714281807
transform 1 0 588 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1592
timestamp 1714281807
transform 1 0 1276 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1593
timestamp 1714281807
transform 1 0 1276 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1594
timestamp 1714281807
transform 1 0 1156 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1595
timestamp 1714281807
transform 1 0 1028 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1596
timestamp 1714281807
transform 1 0 948 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1597
timestamp 1714281807
transform 1 0 1308 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1598
timestamp 1714281807
transform 1 0 1284 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1599
timestamp 1714281807
transform 1 0 1076 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1600
timestamp 1714281807
transform 1 0 1004 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1601
timestamp 1714281807
transform 1 0 1004 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1602
timestamp 1714281807
transform 1 0 1284 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1603
timestamp 1714281807
transform 1 0 1220 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1604
timestamp 1714281807
transform 1 0 1164 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1605
timestamp 1714281807
transform 1 0 1164 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1606
timestamp 1714281807
transform 1 0 1156 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1607
timestamp 1714281807
transform 1 0 1348 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1608
timestamp 1714281807
transform 1 0 1348 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1609
timestamp 1714281807
transform 1 0 1316 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1610
timestamp 1714281807
transform 1 0 1100 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1611
timestamp 1714281807
transform 1 0 1100 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1612
timestamp 1714281807
transform 1 0 500 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1613
timestamp 1714281807
transform 1 0 484 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1614
timestamp 1714281807
transform 1 0 476 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1615
timestamp 1714281807
transform 1 0 484 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1616
timestamp 1714281807
transform 1 0 468 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1617
timestamp 1714281807
transform 1 0 420 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1618
timestamp 1714281807
transform 1 0 420 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1619
timestamp 1714281807
transform 1 0 1756 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1620
timestamp 1714281807
transform 1 0 1740 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1621
timestamp 1714281807
transform 1 0 1676 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1622
timestamp 1714281807
transform 1 0 1564 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1623
timestamp 1714281807
transform 1 0 1564 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1624
timestamp 1714281807
transform 1 0 1636 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1625
timestamp 1714281807
transform 1 0 1612 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1626
timestamp 1714281807
transform 1 0 1596 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1627
timestamp 1714281807
transform 1 0 1548 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1628
timestamp 1714281807
transform 1 0 1828 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1629
timestamp 1714281807
transform 1 0 1828 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1630
timestamp 1714281807
transform 1 0 1700 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1631
timestamp 1714281807
transform 1 0 1700 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1632
timestamp 1714281807
transform 1 0 1612 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1633
timestamp 1714281807
transform 1 0 1596 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1634
timestamp 1714281807
transform 1 0 1828 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1635
timestamp 1714281807
transform 1 0 1828 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1636
timestamp 1714281807
transform 1 0 1796 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1637
timestamp 1714281807
transform 1 0 1764 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1638
timestamp 1714281807
transform 1 0 1380 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1639
timestamp 1714281807
transform 1 0 1356 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1640
timestamp 1714281807
transform 1 0 1156 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1641
timestamp 1714281807
transform 1 0 1092 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1642
timestamp 1714281807
transform 1 0 1092 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1643
timestamp 1714281807
transform 1 0 1092 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1644
timestamp 1714281807
transform 1 0 1212 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1645
timestamp 1714281807
transform 1 0 1084 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1646
timestamp 1714281807
transform 1 0 1084 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1647
timestamp 1714281807
transform 1 0 1220 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1648
timestamp 1714281807
transform 1 0 1220 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1649
timestamp 1714281807
transform 1 0 1220 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1650
timestamp 1714281807
transform 1 0 1204 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1651
timestamp 1714281807
transform 1 0 1316 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1652
timestamp 1714281807
transform 1 0 1180 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1653
timestamp 1714281807
transform 1 0 1076 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1654
timestamp 1714281807
transform 1 0 1044 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1655
timestamp 1714281807
transform 1 0 1100 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1656
timestamp 1714281807
transform 1 0 1060 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1657
timestamp 1714281807
transform 1 0 1052 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1658
timestamp 1714281807
transform 1 0 1380 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1659
timestamp 1714281807
transform 1 0 1380 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1660
timestamp 1714281807
transform 1 0 1372 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1661
timestamp 1714281807
transform 1 0 1332 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1662
timestamp 1714281807
transform 1 0 1764 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1663
timestamp 1714281807
transform 1 0 1732 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1664
timestamp 1714281807
transform 1 0 1732 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1665
timestamp 1714281807
transform 1 0 1676 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1666
timestamp 1714281807
transform 1 0 1548 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1667
timestamp 1714281807
transform 1 0 1540 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1668
timestamp 1714281807
transform 1 0 1500 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1669
timestamp 1714281807
transform 1 0 1500 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1670
timestamp 1714281807
transform 1 0 1876 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1671
timestamp 1714281807
transform 1 0 1860 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1672
timestamp 1714281807
transform 1 0 1820 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1673
timestamp 1714281807
transform 1 0 1820 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1674
timestamp 1714281807
transform 1 0 1788 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1675
timestamp 1714281807
transform 1 0 2132 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1676
timestamp 1714281807
transform 1 0 2084 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1677
timestamp 1714281807
transform 1 0 2036 0 1 295
box -2 -2 2 2
use M2_M1  M2_M1_1678
timestamp 1714281807
transform 1 0 2036 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1679
timestamp 1714281807
transform 1 0 2100 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1680
timestamp 1714281807
transform 1 0 2100 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1681
timestamp 1714281807
transform 1 0 2084 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1682
timestamp 1714281807
transform 1 0 1972 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1683
timestamp 1714281807
transform 1 0 2276 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1684
timestamp 1714281807
transform 1 0 2276 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1685
timestamp 1714281807
transform 1 0 2228 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1686
timestamp 1714281807
transform 1 0 2220 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1687
timestamp 1714281807
transform 1 0 2636 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1688
timestamp 1714281807
transform 1 0 2604 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1689
timestamp 1714281807
transform 1 0 2572 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1690
timestamp 1714281807
transform 1 0 2572 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1691
timestamp 1714281807
transform 1 0 2444 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1692
timestamp 1714281807
transform 1 0 2444 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1693
timestamp 1714281807
transform 1 0 2428 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1694
timestamp 1714281807
transform 1 0 2404 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1695
timestamp 1714281807
transform 1 0 2404 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_1696
timestamp 1714281807
transform 1 0 2732 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1697
timestamp 1714281807
transform 1 0 2700 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_1698
timestamp 1714281807
transform 1 0 2332 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_1699
timestamp 1714281807
transform 1 0 2028 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_1700
timestamp 1714281807
transform 1 0 1956 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1701
timestamp 1714281807
transform 1 0 2020 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1702
timestamp 1714281807
transform 1 0 2020 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1703
timestamp 1714281807
transform 1 0 1972 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1704
timestamp 1714281807
transform 1 0 1940 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1705
timestamp 1714281807
transform 1 0 1940 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1706
timestamp 1714281807
transform 1 0 1804 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_1707
timestamp 1714281807
transform 1 0 1804 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_1708
timestamp 1714281807
transform 1 0 1700 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1709
timestamp 1714281807
transform 1 0 1564 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1710
timestamp 1714281807
transform 1 0 1436 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_1711
timestamp 1714281807
transform 1 0 1500 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1712
timestamp 1714281807
transform 1 0 1436 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1713
timestamp 1714281807
transform 1 0 1436 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1714
timestamp 1714281807
transform 1 0 1260 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_1715
timestamp 1714281807
transform 1 0 684 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1716
timestamp 1714281807
transform 1 0 676 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_1717
timestamp 1714281807
transform 1 0 660 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1718
timestamp 1714281807
transform 1 0 660 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1719
timestamp 1714281807
transform 1 0 700 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1720
timestamp 1714281807
transform 1 0 676 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1721
timestamp 1714281807
transform 1 0 868 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_1722
timestamp 1714281807
transform 1 0 780 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1723
timestamp 1714281807
transform 1 0 1844 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1724
timestamp 1714281807
transform 1 0 1812 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1725
timestamp 1714281807
transform 1 0 1668 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1726
timestamp 1714281807
transform 1 0 2068 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1727
timestamp 1714281807
transform 1 0 2068 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1728
timestamp 1714281807
transform 1 0 2012 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1729
timestamp 1714281807
transform 1 0 2012 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1730
timestamp 1714281807
transform 1 0 1964 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1731
timestamp 1714281807
transform 1 0 1908 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1732
timestamp 1714281807
transform 1 0 1788 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1733
timestamp 1714281807
transform 1 0 1788 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_1734
timestamp 1714281807
transform 1 0 1732 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1735
timestamp 1714281807
transform 1 0 1732 0 1 2045
box -2 -2 2 2
use M2_M1  M2_M1_1736
timestamp 1714281807
transform 1 0 1724 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1737
timestamp 1714281807
transform 1 0 1852 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1738
timestamp 1714281807
transform 1 0 1724 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1739
timestamp 1714281807
transform 1 0 1724 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1740
timestamp 1714281807
transform 1 0 1940 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1741
timestamp 1714281807
transform 1 0 1820 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1742
timestamp 1714281807
transform 1 0 1716 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1743
timestamp 1714281807
transform 1 0 572 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1744
timestamp 1714281807
transform 1 0 540 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1745
timestamp 1714281807
transform 1 0 428 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1746
timestamp 1714281807
transform 1 0 396 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1747
timestamp 1714281807
transform 1 0 1124 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1748
timestamp 1714281807
transform 1 0 1084 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1749
timestamp 1714281807
transform 1 0 1180 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1750
timestamp 1714281807
transform 1 0 1068 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1751
timestamp 1714281807
transform 1 0 772 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1752
timestamp 1714281807
transform 1 0 676 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1753
timestamp 1714281807
transform 1 0 676 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1754
timestamp 1714281807
transform 1 0 652 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1755
timestamp 1714281807
transform 1 0 652 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1756
timestamp 1714281807
transform 1 0 748 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1757
timestamp 1714281807
transform 1 0 740 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1758
timestamp 1714281807
transform 1 0 644 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1759
timestamp 1714281807
transform 1 0 636 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1760
timestamp 1714281807
transform 1 0 636 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1761
timestamp 1714281807
transform 1 0 1132 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1762
timestamp 1714281807
transform 1 0 796 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1763
timestamp 1714281807
transform 1 0 1220 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1764
timestamp 1714281807
transform 1 0 796 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1765
timestamp 1714281807
transform 1 0 636 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1766
timestamp 1714281807
transform 1 0 604 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1767
timestamp 1714281807
transform 1 0 1028 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1768
timestamp 1714281807
transform 1 0 756 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1769
timestamp 1714281807
transform 1 0 1052 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1770
timestamp 1714281807
transform 1 0 788 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1771
timestamp 1714281807
transform 1 0 572 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1772
timestamp 1714281807
transform 1 0 548 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1773
timestamp 1714281807
transform 1 0 1396 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1774
timestamp 1714281807
transform 1 0 1228 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1775
timestamp 1714281807
transform 1 0 1308 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1776
timestamp 1714281807
transform 1 0 1260 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1777
timestamp 1714281807
transform 1 0 1172 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1778
timestamp 1714281807
transform 1 0 1172 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_1779
timestamp 1714281807
transform 1 0 1156 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1780
timestamp 1714281807
transform 1 0 1388 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1781
timestamp 1714281807
transform 1 0 1372 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1782
timestamp 1714281807
transform 1 0 1300 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1783
timestamp 1714281807
transform 1 0 1260 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1784
timestamp 1714281807
transform 1 0 1148 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1785
timestamp 1714281807
transform 1 0 1124 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1786
timestamp 1714281807
transform 1 0 1124 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1787
timestamp 1714281807
transform 1 0 1388 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1788
timestamp 1714281807
transform 1 0 1348 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1789
timestamp 1714281807
transform 1 0 1308 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1790
timestamp 1714281807
transform 1 0 1268 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1791
timestamp 1714281807
transform 1 0 932 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1792
timestamp 1714281807
transform 1 0 828 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1793
timestamp 1714281807
transform 1 0 748 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1794
timestamp 1714281807
transform 1 0 724 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1795
timestamp 1714281807
transform 1 0 1012 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1796
timestamp 1714281807
transform 1 0 964 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1797
timestamp 1714281807
transform 1 0 964 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1798
timestamp 1714281807
transform 1 0 940 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1799
timestamp 1714281807
transform 1 0 908 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1800
timestamp 1714281807
transform 1 0 900 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1801
timestamp 1714281807
transform 1 0 1004 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1802
timestamp 1714281807
transform 1 0 1004 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_1803
timestamp 1714281807
transform 1 0 996 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1804
timestamp 1714281807
transform 1 0 956 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_1805
timestamp 1714281807
transform 1 0 852 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1806
timestamp 1714281807
transform 1 0 748 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1807
timestamp 1714281807
transform 1 0 988 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_1808
timestamp 1714281807
transform 1 0 964 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1809
timestamp 1714281807
transform 1 0 956 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1810
timestamp 1714281807
transform 1 0 796 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_1811
timestamp 1714281807
transform 1 0 660 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1812
timestamp 1714281807
transform 1 0 652 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_1813
timestamp 1714281807
transform 1 0 652 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1814
timestamp 1714281807
transform 1 0 820 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1815
timestamp 1714281807
transform 1 0 756 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_1816
timestamp 1714281807
transform 1 0 564 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1817
timestamp 1714281807
transform 1 0 564 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1818
timestamp 1714281807
transform 1 0 788 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1819
timestamp 1714281807
transform 1 0 556 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1820
timestamp 1714281807
transform 1 0 468 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1821
timestamp 1714281807
transform 1 0 1444 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1822
timestamp 1714281807
transform 1 0 1260 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1823
timestamp 1714281807
transform 1 0 1004 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1824
timestamp 1714281807
transform 1 0 1492 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1825
timestamp 1714281807
transform 1 0 1492 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_1826
timestamp 1714281807
transform 1 0 2228 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1827
timestamp 1714281807
transform 1 0 1468 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1828
timestamp 1714281807
transform 1 0 2236 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1829
timestamp 1714281807
transform 1 0 2204 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1830
timestamp 1714281807
transform 1 0 2212 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1831
timestamp 1714281807
transform 1 0 2212 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1832
timestamp 1714281807
transform 1 0 2380 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1833
timestamp 1714281807
transform 1 0 2220 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_1834
timestamp 1714281807
transform 1 0 2404 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1835
timestamp 1714281807
transform 1 0 2356 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1836
timestamp 1714281807
transform 1 0 2468 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1837
timestamp 1714281807
transform 1 0 2364 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1838
timestamp 1714281807
transform 1 0 2460 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_1839
timestamp 1714281807
transform 1 0 2460 0 1 1245
box -2 -2 2 2
use M2_M1  M2_M1_1840
timestamp 1714281807
transform 1 0 2772 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_1841
timestamp 1714281807
transform 1 0 2540 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1842
timestamp 1714281807
transform 1 0 2876 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1843
timestamp 1714281807
transform 1 0 2756 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_1844
timestamp 1714281807
transform 1 0 2820 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1845
timestamp 1714281807
transform 1 0 2756 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1846
timestamp 1714281807
transform 1 0 2428 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_1847
timestamp 1714281807
transform 1 0 2412 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1848
timestamp 1714281807
transform 1 0 2468 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1849
timestamp 1714281807
transform 1 0 2444 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_1850
timestamp 1714281807
transform 1 0 2412 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_1851
timestamp 1714281807
transform 1 0 1612 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_1852
timestamp 1714281807
transform 1 0 2652 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_1853
timestamp 1714281807
transform 1 0 2500 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1854
timestamp 1714281807
transform 1 0 2876 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1855
timestamp 1714281807
transform 1 0 2628 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_1856
timestamp 1714281807
transform 1 0 2660 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1857
timestamp 1714281807
transform 1 0 2636 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1858
timestamp 1714281807
transform 1 0 2636 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1859
timestamp 1714281807
transform 1 0 2636 0 1 2635
box -2 -2 2 2
use M2_M1  M2_M1_1860
timestamp 1714281807
transform 1 0 1604 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1861
timestamp 1714281807
transform 1 0 1580 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1862
timestamp 1714281807
transform 1 0 1564 0 1 2705
box -2 -2 2 2
use M2_M1  M2_M1_1863
timestamp 1714281807
transform 1 0 1556 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1864
timestamp 1714281807
transform 1 0 2140 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_1865
timestamp 1714281807
transform 1 0 2092 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_1866
timestamp 1714281807
transform 1 0 2204 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_1867
timestamp 1714281807
transform 1 0 2204 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1868
timestamp 1714281807
transform 1 0 2372 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1869
timestamp 1714281807
transform 1 0 2180 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_1870
timestamp 1714281807
transform 1 0 2244 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1871
timestamp 1714281807
transform 1 0 2188 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1872
timestamp 1714281807
transform 1 0 2028 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_1873
timestamp 1714281807
transform 1 0 2020 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1874
timestamp 1714281807
transform 1 0 2028 0 1 2635
box -2 -2 2 2
use M2_M1  M2_M1_1875
timestamp 1714281807
transform 1 0 1908 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1876
timestamp 1714281807
transform 1 0 2044 0 1 2635
box -2 -2 2 2
use M2_M1  M2_M1_1877
timestamp 1714281807
transform 1 0 1876 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1878
timestamp 1714281807
transform 1 0 2628 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1879
timestamp 1714281807
transform 1 0 2292 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_1880
timestamp 1714281807
transform 1 0 2308 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1881
timestamp 1714281807
transform 1 0 2308 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1882
timestamp 1714281807
transform 1 0 2268 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1883
timestamp 1714281807
transform 1 0 2268 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1884
timestamp 1714281807
transform 1 0 2364 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1885
timestamp 1714281807
transform 1 0 2292 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1886
timestamp 1714281807
transform 1 0 2356 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1887
timestamp 1714281807
transform 1 0 2300 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_1888
timestamp 1714281807
transform 1 0 2660 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1889
timestamp 1714281807
transform 1 0 2612 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1890
timestamp 1714281807
transform 1 0 2652 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1891
timestamp 1714281807
transform 1 0 2612 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1892
timestamp 1714281807
transform 1 0 2700 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1893
timestamp 1714281807
transform 1 0 2620 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_1894
timestamp 1714281807
transform 1 0 1460 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_1895
timestamp 1714281807
transform 1 0 1380 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1896
timestamp 1714281807
transform 1 0 1612 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1897
timestamp 1714281807
transform 1 0 1476 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1898
timestamp 1714281807
transform 1 0 1836 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1899
timestamp 1714281807
transform 1 0 1484 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_1900
timestamp 1714281807
transform 1 0 2388 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1901
timestamp 1714281807
transform 1 0 1796 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1902
timestamp 1714281807
transform 1 0 1804 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1903
timestamp 1714281807
transform 1 0 1788 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_1904
timestamp 1714281807
transform 1 0 1732 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_1905
timestamp 1714281807
transform 1 0 1668 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1906
timestamp 1714281807
transform 1 0 1948 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1907
timestamp 1714281807
transform 1 0 1788 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1908
timestamp 1714281807
transform 1 0 1996 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1909
timestamp 1714281807
transform 1 0 1924 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1910
timestamp 1714281807
transform 1 0 1932 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1911
timestamp 1714281807
transform 1 0 1788 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1912
timestamp 1714281807
transform 1 0 2268 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1913
timestamp 1714281807
transform 1 0 1940 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_1914
timestamp 1714281807
transform 1 0 1596 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1915
timestamp 1714281807
transform 1 0 1572 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1916
timestamp 1714281807
transform 1 0 1596 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1917
timestamp 1714281807
transform 1 0 1412 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1918
timestamp 1714281807
transform 1 0 1812 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1919
timestamp 1714281807
transform 1 0 1612 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_1920
timestamp 1714281807
transform 1 0 2396 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1921
timestamp 1714281807
transform 1 0 2380 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_1922
timestamp 1714281807
transform 1 0 2676 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1923
timestamp 1714281807
transform 1 0 2452 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1924
timestamp 1714281807
transform 1 0 2684 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1925
timestamp 1714281807
transform 1 0 2660 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1926
timestamp 1714281807
transform 1 0 2932 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1927
timestamp 1714281807
transform 1 0 2668 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_1928
timestamp 1714281807
transform 1 0 2436 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1929
timestamp 1714281807
transform 1 0 2380 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1930
timestamp 1714281807
transform 1 0 2380 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1931
timestamp 1714281807
transform 1 0 2188 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1932
timestamp 1714281807
transform 1 0 2668 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1933
timestamp 1714281807
transform 1 0 2388 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_1934
timestamp 1714281807
transform 1 0 1628 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_1935
timestamp 1714281807
transform 1 0 1628 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_1936
timestamp 1714281807
transform 1 0 1716 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_1937
timestamp 1714281807
transform 1 0 1684 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_1938
timestamp 1714281807
transform 1 0 1820 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1939
timestamp 1714281807
transform 1 0 1700 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_1940
timestamp 1714281807
transform 1 0 1708 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1941
timestamp 1714281807
transform 1 0 1700 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1942
timestamp 1714281807
transform 1 0 1652 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_1943
timestamp 1714281807
transform 1 0 1412 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1944
timestamp 1714281807
transform 1 0 1636 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1945
timestamp 1714281807
transform 1 0 1564 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_1946
timestamp 1714281807
transform 1 0 1596 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1947
timestamp 1714281807
transform 1 0 1572 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_1948
timestamp 1714281807
transform 1 0 1860 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1949
timestamp 1714281807
transform 1 0 1636 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_1950
timestamp 1714281807
transform 1 0 1700 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1951
timestamp 1714281807
transform 1 0 1676 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1952
timestamp 1714281807
transform 1 0 1396 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1953
timestamp 1714281807
transform 1 0 1236 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_1954
timestamp 1714281807
transform 1 0 1188 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_1955
timestamp 1714281807
transform 1 0 1188 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1956
timestamp 1714281807
transform 1 0 1356 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1957
timestamp 1714281807
transform 1 0 1204 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_1958
timestamp 1714281807
transform 1 0 1628 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1959
timestamp 1714281807
transform 1 0 1324 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1960
timestamp 1714281807
transform 1 0 1300 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_1961
timestamp 1714281807
transform 1 0 1252 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1962
timestamp 1714281807
transform 1 0 1420 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1963
timestamp 1714281807
transform 1 0 964 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_1964
timestamp 1714281807
transform 1 0 940 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1965
timestamp 1714281807
transform 1 0 836 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_1966
timestamp 1714281807
transform 1 0 724 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_1967
timestamp 1714281807
transform 1 0 644 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1968
timestamp 1714281807
transform 1 0 892 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_1969
timestamp 1714281807
transform 1 0 852 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1970
timestamp 1714281807
transform 1 0 2564 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1971
timestamp 1714281807
transform 1 0 2564 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1972
timestamp 1714281807
transform 1 0 2516 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1973
timestamp 1714281807
transform 1 0 2492 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1974
timestamp 1714281807
transform 1 0 2484 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1975
timestamp 1714281807
transform 1 0 2356 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1976
timestamp 1714281807
transform 1 0 2300 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1977
timestamp 1714281807
transform 1 0 2300 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1978
timestamp 1714281807
transform 1 0 1508 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1979
timestamp 1714281807
transform 1 0 2516 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1980
timestamp 1714281807
transform 1 0 2476 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1981
timestamp 1714281807
transform 1 0 2500 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1982
timestamp 1714281807
transform 1 0 2404 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1983
timestamp 1714281807
transform 1 0 2372 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1984
timestamp 1714281807
transform 1 0 2268 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1985
timestamp 1714281807
transform 1 0 2596 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1986
timestamp 1714281807
transform 1 0 2548 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1987
timestamp 1714281807
transform 1 0 2316 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1988
timestamp 1714281807
transform 1 0 2284 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1989
timestamp 1714281807
transform 1 0 1436 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1990
timestamp 1714281807
transform 1 0 1140 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1991
timestamp 1714281807
transform 1 0 1236 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1992
timestamp 1714281807
transform 1 0 1212 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1993
timestamp 1714281807
transform 1 0 1044 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1994
timestamp 1714281807
transform 1 0 1172 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1995
timestamp 1714281807
transform 1 0 1084 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1996
timestamp 1714281807
transform 1 0 1084 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1997
timestamp 1714281807
transform 1 0 1076 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1998
timestamp 1714281807
transform 1 0 1004 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1999
timestamp 1714281807
transform 1 0 1148 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2000
timestamp 1714281807
transform 1 0 748 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2001
timestamp 1714281807
transform 1 0 476 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2002
timestamp 1714281807
transform 1 0 2108 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2003
timestamp 1714281807
transform 1 0 2108 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2004
timestamp 1714281807
transform 1 0 2052 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2005
timestamp 1714281807
transform 1 0 2044 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2006
timestamp 1714281807
transform 1 0 1940 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2007
timestamp 1714281807
transform 1 0 1908 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2008
timestamp 1714281807
transform 1 0 1868 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2009
timestamp 1714281807
transform 1 0 1140 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2010
timestamp 1714281807
transform 1 0 2124 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2011
timestamp 1714281807
transform 1 0 2012 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2012
timestamp 1714281807
transform 1 0 2044 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2013
timestamp 1714281807
transform 1 0 1956 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2014
timestamp 1714281807
transform 1 0 1876 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2015
timestamp 1714281807
transform 1 0 2100 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2016
timestamp 1714281807
transform 1 0 2092 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2017
timestamp 1714281807
transform 1 0 1892 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2018
timestamp 1714281807
transform 1 0 1884 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2019
timestamp 1714281807
transform 1 0 1108 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2020
timestamp 1714281807
transform 1 0 1092 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2021
timestamp 1714281807
transform 1 0 1036 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2022
timestamp 1714281807
transform 1 0 620 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2023
timestamp 1714281807
transform 1 0 324 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2024
timestamp 1714281807
transform 1 0 1716 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2025
timestamp 1714281807
transform 1 0 1660 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2026
timestamp 1714281807
transform 1 0 1556 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2027
timestamp 1714281807
transform 1 0 1476 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2028
timestamp 1714281807
transform 1 0 1476 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2029
timestamp 1714281807
transform 1 0 1436 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2030
timestamp 1714281807
transform 1 0 1436 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2031
timestamp 1714281807
transform 1 0 1420 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2032
timestamp 1714281807
transform 1 0 1244 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2033
timestamp 1714281807
transform 1 0 1548 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2034
timestamp 1714281807
transform 1 0 1524 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2035
timestamp 1714281807
transform 1 0 1692 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2036
timestamp 1714281807
transform 1 0 1492 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2037
timestamp 1714281807
transform 1 0 1412 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2038
timestamp 1714281807
transform 1 0 1724 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2039
timestamp 1714281807
transform 1 0 1708 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2040
timestamp 1714281807
transform 1 0 1444 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2041
timestamp 1714281807
transform 1 0 1428 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2042
timestamp 1714281807
transform 1 0 1180 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2043
timestamp 1714281807
transform 1 0 1164 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2044
timestamp 1714281807
transform 1 0 1004 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2045
timestamp 1714281807
transform 1 0 708 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2046
timestamp 1714281807
transform 1 0 260 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2047
timestamp 1714281807
transform 1 0 1292 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2048
timestamp 1714281807
transform 1 0 1276 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2049
timestamp 1714281807
transform 1 0 1212 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2050
timestamp 1714281807
transform 1 0 1212 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2051
timestamp 1714281807
transform 1 0 1156 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2052
timestamp 1714281807
transform 1 0 1076 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2053
timestamp 1714281807
transform 1 0 1068 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2054
timestamp 1714281807
transform 1 0 1060 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2055
timestamp 1714281807
transform 1 0 1148 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2056
timestamp 1714281807
transform 1 0 1124 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2057
timestamp 1714281807
transform 1 0 1228 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2058
timestamp 1714281807
transform 1 0 1132 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2059
timestamp 1714281807
transform 1 0 1132 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_2060
timestamp 1714281807
transform 1 0 1196 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2061
timestamp 1714281807
transform 1 0 1172 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2062
timestamp 1714281807
transform 1 0 1292 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2063
timestamp 1714281807
transform 1 0 1284 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2064
timestamp 1714281807
transform 1 0 1052 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2065
timestamp 1714281807
transform 1 0 1036 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2066
timestamp 1714281807
transform 1 0 1148 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2067
timestamp 1714281807
transform 1 0 1100 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2068
timestamp 1714281807
transform 1 0 996 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2069
timestamp 1714281807
transform 1 0 964 0 1 1585
box -2 -2 2 2
use M2_M1  M2_M1_2070
timestamp 1714281807
transform 1 0 964 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_2071
timestamp 1714281807
transform 1 0 964 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2072
timestamp 1714281807
transform 1 0 764 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2073
timestamp 1714281807
transform 1 0 508 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2074
timestamp 1714281807
transform 1 0 252 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2075
timestamp 1714281807
transform 1 0 1268 0 1 985
box -2 -2 2 2
use M2_M1  M2_M1_2076
timestamp 1714281807
transform 1 0 1220 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2077
timestamp 1714281807
transform 1 0 1204 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2078
timestamp 1714281807
transform 1 0 1204 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2079
timestamp 1714281807
transform 1 0 1116 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2080
timestamp 1714281807
transform 1 0 1116 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2081
timestamp 1714281807
transform 1 0 1100 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2082
timestamp 1714281807
transform 1 0 1100 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2083
timestamp 1714281807
transform 1 0 1196 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2084
timestamp 1714281807
transform 1 0 1172 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2085
timestamp 1714281807
transform 1 0 1236 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2086
timestamp 1714281807
transform 1 0 1220 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2087
timestamp 1714281807
transform 1 0 1172 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2088
timestamp 1714281807
transform 1 0 1172 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2089
timestamp 1714281807
transform 1 0 1188 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2090
timestamp 1714281807
transform 1 0 1164 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2091
timestamp 1714281807
transform 1 0 1244 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2092
timestamp 1714281807
transform 1 0 1220 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2093
timestamp 1714281807
transform 1 0 1092 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_2094
timestamp 1714281807
transform 1 0 1012 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2095
timestamp 1714281807
transform 1 0 724 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2096
timestamp 1714281807
transform 1 0 564 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2097
timestamp 1714281807
transform 1 0 404 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2098
timestamp 1714281807
transform 1 0 1852 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2099
timestamp 1714281807
transform 1 0 1836 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2100
timestamp 1714281807
transform 1 0 1836 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2101
timestamp 1714281807
transform 1 0 1788 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2102
timestamp 1714281807
transform 1 0 1756 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2103
timestamp 1714281807
transform 1 0 1756 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2104
timestamp 1714281807
transform 1 0 1620 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2105
timestamp 1714281807
transform 1 0 1532 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2106
timestamp 1714281807
transform 1 0 1852 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2107
timestamp 1714281807
transform 1 0 1844 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2108
timestamp 1714281807
transform 1 0 1772 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2109
timestamp 1714281807
transform 1 0 1764 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2110
timestamp 1714281807
transform 1 0 1692 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2111
timestamp 1714281807
transform 1 0 1708 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2112
timestamp 1714281807
transform 1 0 1684 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2113
timestamp 1714281807
transform 1 0 1860 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_2114
timestamp 1714281807
transform 1 0 1780 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2115
timestamp 1714281807
transform 1 0 1388 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2116
timestamp 1714281807
transform 1 0 1116 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2117
timestamp 1714281807
transform 1 0 764 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2118
timestamp 1714281807
transform 1 0 620 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2119
timestamp 1714281807
transform 1 0 444 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2120
timestamp 1714281807
transform 1 0 1756 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2121
timestamp 1714281807
transform 1 0 1692 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2122
timestamp 1714281807
transform 1 0 1684 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2123
timestamp 1714281807
transform 1 0 1676 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2124
timestamp 1714281807
transform 1 0 1572 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2125
timestamp 1714281807
transform 1 0 1516 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2126
timestamp 1714281807
transform 1 0 1508 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2127
timestamp 1714281807
transform 1 0 1660 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2128
timestamp 1714281807
transform 1 0 1636 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2129
timestamp 1714281807
transform 1 0 1700 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2130
timestamp 1714281807
transform 1 0 1652 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2131
timestamp 1714281807
transform 1 0 1644 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2132
timestamp 1714281807
transform 1 0 1668 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2133
timestamp 1714281807
transform 1 0 1644 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2134
timestamp 1714281807
transform 1 0 1764 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2135
timestamp 1714281807
transform 1 0 1748 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2136
timestamp 1714281807
transform 1 0 1460 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2137
timestamp 1714281807
transform 1 0 1204 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2138
timestamp 1714281807
transform 1 0 748 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2139
timestamp 1714281807
transform 1 0 652 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2140
timestamp 1714281807
transform 1 0 588 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2141
timestamp 1714281807
transform 1 0 924 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2142
timestamp 1714281807
transform 1 0 924 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2143
timestamp 1714281807
transform 1 0 2420 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2144
timestamp 1714281807
transform 1 0 2380 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2145
timestamp 1714281807
transform 1 0 2380 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2146
timestamp 1714281807
transform 1 0 2340 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2147
timestamp 1714281807
transform 1 0 2260 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2148
timestamp 1714281807
transform 1 0 2236 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2149
timestamp 1714281807
transform 1 0 1564 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2150
timestamp 1714281807
transform 1 0 2396 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2151
timestamp 1714281807
transform 1 0 2252 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2152
timestamp 1714281807
transform 1 0 2292 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2153
timestamp 1714281807
transform 1 0 2292 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2154
timestamp 1714281807
transform 1 0 2252 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2155
timestamp 1714281807
transform 1 0 2236 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2156
timestamp 1714281807
transform 1 0 2444 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2157
timestamp 1714281807
transform 1 0 2340 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2158
timestamp 1714281807
transform 1 0 2436 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2159
timestamp 1714281807
transform 1 0 2332 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2160
timestamp 1714281807
transform 1 0 1484 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2161
timestamp 1714281807
transform 1 0 1284 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2162
timestamp 1714281807
transform 1 0 1316 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2163
timestamp 1714281807
transform 1 0 1316 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2164
timestamp 1714281807
transform 1 0 1252 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2165
timestamp 1714281807
transform 1 0 1252 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2166
timestamp 1714281807
transform 1 0 1020 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2167
timestamp 1714281807
transform 1 0 1196 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2168
timestamp 1714281807
transform 1 0 1116 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2169
timestamp 1714281807
transform 1 0 1092 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2170
timestamp 1714281807
transform 1 0 2860 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2171
timestamp 1714281807
transform 1 0 2828 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2172
timestamp 1714281807
transform 1 0 2772 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2173
timestamp 1714281807
transform 1 0 2764 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2174
timestamp 1714281807
transform 1 0 2756 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2175
timestamp 1714281807
transform 1 0 2692 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2176
timestamp 1714281807
transform 1 0 1492 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2177
timestamp 1714281807
transform 1 0 2868 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2178
timestamp 1714281807
transform 1 0 2764 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2179
timestamp 1714281807
transform 1 0 2788 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2180
timestamp 1714281807
transform 1 0 2724 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2181
timestamp 1714281807
transform 1 0 2724 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2182
timestamp 1714281807
transform 1 0 2780 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_2183
timestamp 1714281807
transform 1 0 2740 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2184
timestamp 1714281807
transform 1 0 2908 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2185
timestamp 1714281807
transform 1 0 2820 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2186
timestamp 1714281807
transform 1 0 1436 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2187
timestamp 1714281807
transform 1 0 1372 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2188
timestamp 1714281807
transform 1 0 1316 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2189
timestamp 1714281807
transform 1 0 1156 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2190
timestamp 1714281807
transform 1 0 1140 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_2191
timestamp 1714281807
transform 1 0 2428 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2192
timestamp 1714281807
transform 1 0 2396 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_2193
timestamp 1714281807
transform 1 0 2308 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_2194
timestamp 1714281807
transform 1 0 2252 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2195
timestamp 1714281807
transform 1 0 2228 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2196
timestamp 1714281807
transform 1 0 2124 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_2197
timestamp 1714281807
transform 1 0 2060 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2198
timestamp 1714281807
transform 1 0 1404 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2199
timestamp 1714281807
transform 1 0 2316 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_2200
timestamp 1714281807
transform 1 0 2300 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2201
timestamp 1714281807
transform 1 0 2324 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2202
timestamp 1714281807
transform 1 0 2244 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2203
timestamp 1714281807
transform 1 0 2100 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2204
timestamp 1714281807
transform 1 0 2116 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2205
timestamp 1714281807
transform 1 0 2092 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_2206
timestamp 1714281807
transform 1 0 2444 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_2207
timestamp 1714281807
transform 1 0 2388 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2208
timestamp 1714281807
transform 1 0 1380 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2209
timestamp 1714281807
transform 1 0 1380 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2210
timestamp 1714281807
transform 1 0 1188 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2211
timestamp 1714281807
transform 1 0 1180 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2212
timestamp 1714281807
transform 1 0 1148 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2213
timestamp 1714281807
transform 1 0 1940 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_2214
timestamp 1714281807
transform 1 0 1900 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2215
timestamp 1714281807
transform 1 0 1884 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2216
timestamp 1714281807
transform 1 0 1820 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_2217
timestamp 1714281807
transform 1 0 1756 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2218
timestamp 1714281807
transform 1 0 1740 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_2219
timestamp 1714281807
transform 1 0 1652 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2220
timestamp 1714281807
transform 1 0 1388 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2221
timestamp 1714281807
transform 1 0 1900 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_2222
timestamp 1714281807
transform 1 0 1812 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2223
timestamp 1714281807
transform 1 0 1916 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2224
timestamp 1714281807
transform 1 0 1756 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2225
timestamp 1714281807
transform 1 0 1716 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2226
timestamp 1714281807
transform 1 0 1788 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_2227
timestamp 1714281807
transform 1 0 1732 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2228
timestamp 1714281807
transform 1 0 1988 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_2229
timestamp 1714281807
transform 1 0 1932 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2230
timestamp 1714281807
transform 1 0 1324 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2231
timestamp 1714281807
transform 1 0 1292 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2232
timestamp 1714281807
transform 1 0 1244 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_2233
timestamp 1714281807
transform 1 0 1236 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2234
timestamp 1714281807
transform 1 0 1236 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2235
timestamp 1714281807
transform 1 0 988 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2236
timestamp 1714281807
transform 1 0 972 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2237
timestamp 1714281807
transform 1 0 892 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2238
timestamp 1714281807
transform 1 0 2828 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_2239
timestamp 1714281807
transform 1 0 2772 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2240
timestamp 1714281807
transform 1 0 2724 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_2241
timestamp 1714281807
transform 1 0 2692 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2242
timestamp 1714281807
transform 1 0 2580 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2243
timestamp 1714281807
transform 1 0 2532 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_2244
timestamp 1714281807
transform 1 0 2508 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2245
timestamp 1714281807
transform 1 0 1364 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2246
timestamp 1714281807
transform 1 0 2756 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_2247
timestamp 1714281807
transform 1 0 2716 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2248
timestamp 1714281807
transform 1 0 2740 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2249
timestamp 1714281807
transform 1 0 2668 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2250
timestamp 1714281807
transform 1 0 2596 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2251
timestamp 1714281807
transform 1 0 2508 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2252
timestamp 1714281807
transform 1 0 2532 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_2253
timestamp 1714281807
transform 1 0 2524 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2254
timestamp 1714281807
transform 1 0 2828 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_2255
timestamp 1714281807
transform 1 0 2804 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2256
timestamp 1714281807
transform 1 0 1292 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2257
timestamp 1714281807
transform 1 0 1284 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2258
timestamp 1714281807
transform 1 0 1356 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2259
timestamp 1714281807
transform 1 0 1276 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2260
timestamp 1714281807
transform 1 0 1268 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2261
timestamp 1714281807
transform 1 0 1268 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2262
timestamp 1714281807
transform 1 0 1028 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2263
timestamp 1714281807
transform 1 0 1292 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2264
timestamp 1714281807
transform 1 0 1012 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2265
timestamp 1714281807
transform 1 0 916 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2266
timestamp 1714281807
transform 1 0 1484 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2267
timestamp 1714281807
transform 1 0 1436 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_2268
timestamp 1714281807
transform 1 0 1428 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2269
timestamp 1714281807
transform 1 0 1428 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2270
timestamp 1714281807
transform 1 0 1372 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2271
timestamp 1714281807
transform 1 0 1364 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2272
timestamp 1714281807
transform 1 0 1252 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2273
timestamp 1714281807
transform 1 0 1252 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2274
timestamp 1714281807
transform 1 0 1428 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2275
timestamp 1714281807
transform 1 0 1356 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_2276
timestamp 1714281807
transform 1 0 1428 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2277
timestamp 1714281807
transform 1 0 1380 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2278
timestamp 1714281807
transform 1 0 1380 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2279
timestamp 1714281807
transform 1 0 1476 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_2280
timestamp 1714281807
transform 1 0 1476 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2281
timestamp 1714281807
transform 1 0 1404 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2282
timestamp 1714281807
transform 1 0 1396 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_2283
timestamp 1714281807
transform 1 0 1292 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2284
timestamp 1714281807
transform 1 0 1260 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2285
timestamp 1714281807
transform 1 0 1300 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2286
timestamp 1714281807
transform 1 0 924 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2287
timestamp 1714281807
transform 1 0 796 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2288
timestamp 1714281807
transform 1 0 1012 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2289
timestamp 1714281807
transform 1 0 956 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2290
timestamp 1714281807
transform 1 0 876 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2291
timestamp 1714281807
transform 1 0 436 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2292
timestamp 1714281807
transform 1 0 420 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2293
timestamp 1714281807
transform 1 0 348 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2294
timestamp 1714281807
transform 1 0 2780 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2295
timestamp 1714281807
transform 1 0 2764 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2296
timestamp 1714281807
transform 1 0 2572 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2297
timestamp 1714281807
transform 1 0 2556 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2298
timestamp 1714281807
transform 1 0 1372 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2299
timestamp 1714281807
transform 1 0 2852 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2300
timestamp 1714281807
transform 1 0 2756 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2301
timestamp 1714281807
transform 1 0 2740 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2302
timestamp 1714281807
transform 1 0 2740 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2303
timestamp 1714281807
transform 1 0 2700 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2304
timestamp 1714281807
transform 1 0 2572 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2305
timestamp 1714281807
transform 1 0 2548 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2306
timestamp 1714281807
transform 1 0 2652 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_2307
timestamp 1714281807
transform 1 0 2564 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2308
timestamp 1714281807
transform 1 0 2860 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2309
timestamp 1714281807
transform 1 0 2756 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2310
timestamp 1714281807
transform 1 0 1372 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2311
timestamp 1714281807
transform 1 0 1364 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2312
timestamp 1714281807
transform 1 0 1252 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2313
timestamp 1714281807
transform 1 0 1244 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2314
timestamp 1714281807
transform 1 0 1084 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2315
timestamp 1714281807
transform 1 0 1124 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2316
timestamp 1714281807
transform 1 0 1076 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2317
timestamp 1714281807
transform 1 0 892 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2318
timestamp 1714281807
transform 1 0 492 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2319
timestamp 1714281807
transform 1 0 404 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2320
timestamp 1714281807
transform 1 0 292 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2321
timestamp 1714281807
transform 1 0 2324 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2322
timestamp 1714281807
transform 1 0 2308 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2323
timestamp 1714281807
transform 1 0 2308 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2324
timestamp 1714281807
transform 1 0 2220 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2325
timestamp 1714281807
transform 1 0 2204 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2326
timestamp 1714281807
transform 1 0 2148 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2327
timestamp 1714281807
transform 1 0 1484 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2328
timestamp 1714281807
transform 1 0 2364 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2329
timestamp 1714281807
transform 1 0 2300 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2330
timestamp 1714281807
transform 1 0 2228 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2331
timestamp 1714281807
transform 1 0 2220 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2332
timestamp 1714281807
transform 1 0 2196 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2333
timestamp 1714281807
transform 1 0 2212 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2334
timestamp 1714281807
transform 1 0 2188 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2335
timestamp 1714281807
transform 1 0 2348 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2336
timestamp 1714281807
transform 1 0 2300 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2337
timestamp 1714281807
transform 1 0 1444 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2338
timestamp 1714281807
transform 1 0 1292 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2339
timestamp 1714281807
transform 1 0 1204 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2340
timestamp 1714281807
transform 1 0 980 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2341
timestamp 1714281807
transform 1 0 868 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2342
timestamp 1714281807
transform 1 0 1140 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2343
timestamp 1714281807
transform 1 0 1060 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2344
timestamp 1714281807
transform 1 0 908 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2345
timestamp 1714281807
transform 1 0 548 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2346
timestamp 1714281807
transform 1 0 508 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2347
timestamp 1714281807
transform 1 0 260 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2348
timestamp 1714281807
transform 1 0 900 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2349
timestamp 1714281807
transform 1 0 884 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2350
timestamp 1714281807
transform 1 0 868 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2351
timestamp 1714281807
transform 1 0 2828 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2352
timestamp 1714281807
transform 1 0 2828 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2353
timestamp 1714281807
transform 1 0 2772 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2354
timestamp 1714281807
transform 1 0 2764 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2355
timestamp 1714281807
transform 1 0 2748 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2356
timestamp 1714281807
transform 1 0 2748 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2357
timestamp 1714281807
transform 1 0 2620 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2358
timestamp 1714281807
transform 1 0 1420 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2359
timestamp 1714281807
transform 1 0 2852 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2360
timestamp 1714281807
transform 1 0 2820 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2361
timestamp 1714281807
transform 1 0 2764 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2362
timestamp 1714281807
transform 1 0 2724 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2363
timestamp 1714281807
transform 1 0 2724 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2364
timestamp 1714281807
transform 1 0 2692 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2365
timestamp 1714281807
transform 1 0 2660 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2366
timestamp 1714281807
transform 1 0 940 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_2367
timestamp 1714281807
transform 1 0 940 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2368
timestamp 1714281807
transform 1 0 884 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2369
timestamp 1714281807
transform 1 0 852 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_2370
timestamp 1714281807
transform 1 0 956 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2371
timestamp 1714281807
transform 1 0 948 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2372
timestamp 1714281807
transform 1 0 924 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2373
timestamp 1714281807
transform 1 0 828 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2374
timestamp 1714281807
transform 1 0 828 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2375
timestamp 1714281807
transform 1 0 2764 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2376
timestamp 1714281807
transform 1 0 2740 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2377
timestamp 1714281807
transform 1 0 884 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2378
timestamp 1714281807
transform 1 0 844 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2379
timestamp 1714281807
transform 1 0 844 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2380
timestamp 1714281807
transform 1 0 2860 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2381
timestamp 1714281807
transform 1 0 2764 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2382
timestamp 1714281807
transform 1 0 1388 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2383
timestamp 1714281807
transform 1 0 1236 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2384
timestamp 1714281807
transform 1 0 1244 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2385
timestamp 1714281807
transform 1 0 676 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2386
timestamp 1714281807
transform 1 0 620 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2387
timestamp 1714281807
transform 1 0 1260 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2388
timestamp 1714281807
transform 1 0 1260 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2389
timestamp 1714281807
transform 1 0 1220 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2390
timestamp 1714281807
transform 1 0 1188 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2391
timestamp 1714281807
transform 1 0 860 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2392
timestamp 1714281807
transform 1 0 700 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2393
timestamp 1714281807
transform 1 0 300 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2394
timestamp 1714281807
transform 1 0 268 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2395
timestamp 1714281807
transform 1 0 244 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2396
timestamp 1714281807
transform 1 0 924 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2397
timestamp 1714281807
transform 1 0 924 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2398
timestamp 1714281807
transform 1 0 892 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2399
timestamp 1714281807
transform 1 0 804 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2400
timestamp 1714281807
transform 1 0 492 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2401
timestamp 1714281807
transform 1 0 420 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2402
timestamp 1714281807
transform 1 0 404 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2403
timestamp 1714281807
transform 1 0 836 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2404
timestamp 1714281807
transform 1 0 796 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2405
timestamp 1714281807
transform 1 0 740 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2406
timestamp 1714281807
transform 1 0 436 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2407
timestamp 1714281807
transform 1 0 876 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2408
timestamp 1714281807
transform 1 0 860 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2409
timestamp 1714281807
transform 1 0 1036 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2410
timestamp 1714281807
transform 1 0 860 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2411
timestamp 1714281807
transform 1 0 964 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2412
timestamp 1714281807
transform 1 0 868 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2413
timestamp 1714281807
transform 1 0 948 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2414
timestamp 1714281807
transform 1 0 900 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2415
timestamp 1714281807
transform 1 0 884 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2416
timestamp 1714281807
transform 1 0 868 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2417
timestamp 1714281807
transform 1 0 1108 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2418
timestamp 1714281807
transform 1 0 1036 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2419
timestamp 1714281807
transform 1 0 564 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2420
timestamp 1714281807
transform 1 0 428 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2421
timestamp 1714281807
transform 1 0 532 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2422
timestamp 1714281807
transform 1 0 500 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2423
timestamp 1714281807
transform 1 0 444 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2424
timestamp 1714281807
transform 1 0 428 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2425
timestamp 1714281807
transform 1 0 604 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2426
timestamp 1714281807
transform 1 0 532 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2427
timestamp 1714281807
transform 1 0 300 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2428
timestamp 1714281807
transform 1 0 276 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2429
timestamp 1714281807
transform 1 0 628 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2430
timestamp 1714281807
transform 1 0 628 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2431
timestamp 1714281807
transform 1 0 596 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2432
timestamp 1714281807
transform 1 0 596 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2433
timestamp 1714281807
transform 1 0 548 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2434
timestamp 1714281807
transform 1 0 484 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2435
timestamp 1714281807
transform 1 0 444 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2436
timestamp 1714281807
transform 1 0 716 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2437
timestamp 1714281807
transform 1 0 708 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2438
timestamp 1714281807
transform 1 0 636 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2439
timestamp 1714281807
transform 1 0 620 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2440
timestamp 1714281807
transform 1 0 532 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2441
timestamp 1714281807
transform 1 0 460 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2442
timestamp 1714281807
transform 1 0 692 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2443
timestamp 1714281807
transform 1 0 588 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_2444
timestamp 1714281807
transform 1 0 556 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_2445
timestamp 1714281807
transform 1 0 540 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2446
timestamp 1714281807
transform 1 0 564 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2447
timestamp 1714281807
transform 1 0 532 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2448
timestamp 1714281807
transform 1 0 532 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2449
timestamp 1714281807
transform 1 0 620 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2450
timestamp 1714281807
transform 1 0 556 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2451
timestamp 1714281807
transform 1 0 548 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2452
timestamp 1714281807
transform 1 0 484 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2453
timestamp 1714281807
transform 1 0 2156 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2454
timestamp 1714281807
transform 1 0 2132 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2455
timestamp 1714281807
transform 1 0 2116 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2456
timestamp 1714281807
transform 1 0 2020 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2457
timestamp 1714281807
transform 1 0 2772 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2458
timestamp 1714281807
transform 1 0 2756 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2459
timestamp 1714281807
transform 1 0 2444 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_2460
timestamp 1714281807
transform 1 0 2052 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2461
timestamp 1714281807
transform 1 0 2052 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2462
timestamp 1714281807
transform 1 0 2772 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2463
timestamp 1714281807
transform 1 0 2748 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2464
timestamp 1714281807
transform 1 0 2468 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2465
timestamp 1714281807
transform 1 0 2028 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2466
timestamp 1714281807
transform 1 0 1916 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2467
timestamp 1714281807
transform 1 0 2660 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2468
timestamp 1714281807
transform 1 0 2444 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2469
timestamp 1714281807
transform 1 0 2372 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2470
timestamp 1714281807
transform 1 0 2188 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2471
timestamp 1714281807
transform 1 0 1956 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2472
timestamp 1714281807
transform 1 0 2668 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2473
timestamp 1714281807
transform 1 0 2500 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2474
timestamp 1714281807
transform 1 0 2164 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2475
timestamp 1714281807
transform 1 0 2108 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2476
timestamp 1714281807
transform 1 0 2020 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2477
timestamp 1714281807
transform 1 0 2516 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2478
timestamp 1714281807
transform 1 0 2340 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2479
timestamp 1714281807
transform 1 0 2164 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2480
timestamp 1714281807
transform 1 0 2020 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2481
timestamp 1714281807
transform 1 0 1836 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2482
timestamp 1714281807
transform 1 0 2052 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2483
timestamp 1714281807
transform 1 0 1980 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_2484
timestamp 1714281807
transform 1 0 1948 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2485
timestamp 1714281807
transform 1 0 1444 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_2486
timestamp 1714281807
transform 1 0 1428 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2487
timestamp 1714281807
transform 1 0 2116 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2488
timestamp 1714281807
transform 1 0 1916 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2489
timestamp 1714281807
transform 1 0 1900 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2490
timestamp 1714281807
transform 1 0 1756 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2491
timestamp 1714281807
transform 1 0 1572 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2492
timestamp 1714281807
transform 1 0 2716 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_2493
timestamp 1714281807
transform 1 0 2364 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_2494
timestamp 1714281807
transform 1 0 2028 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2495
timestamp 1714281807
transform 1 0 1780 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2496
timestamp 1714281807
transform 1 0 1500 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2497
timestamp 1714281807
transform 1 0 2620 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_2498
timestamp 1714281807
transform 1 0 2260 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_2499
timestamp 1714281807
transform 1 0 1988 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2500
timestamp 1714281807
transform 1 0 1700 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2501
timestamp 1714281807
transform 1 0 1420 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2502
timestamp 1714281807
transform 1 0 2500 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_2503
timestamp 1714281807
transform 1 0 2140 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_2504
timestamp 1714281807
transform 1 0 1892 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2505
timestamp 1714281807
transform 1 0 1556 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2506
timestamp 1714281807
transform 1 0 1556 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2507
timestamp 1714281807
transform 1 0 2044 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2508
timestamp 1714281807
transform 1 0 2004 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2509
timestamp 1714281807
transform 1 0 1932 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2510
timestamp 1714281807
transform 1 0 1964 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2511
timestamp 1714281807
transform 1 0 1916 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2512
timestamp 1714281807
transform 1 0 1916 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2513
timestamp 1714281807
transform 1 0 1900 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2514
timestamp 1714281807
transform 1 0 2060 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2515
timestamp 1714281807
transform 1 0 2036 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2516
timestamp 1714281807
transform 1 0 1972 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2517
timestamp 1714281807
transform 1 0 1964 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2518
timestamp 1714281807
transform 1 0 1860 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2519
timestamp 1714281807
transform 1 0 1828 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_2520
timestamp 1714281807
transform 1 0 1740 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_2521
timestamp 1714281807
transform 1 0 1980 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2522
timestamp 1714281807
transform 1 0 1972 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2523
timestamp 1714281807
transform 1 0 1924 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2524
timestamp 1714281807
transform 1 0 1884 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2525
timestamp 1714281807
transform 1 0 1820 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2526
timestamp 1714281807
transform 1 0 1804 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_2527
timestamp 1714281807
transform 1 0 1644 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2528
timestamp 1714281807
transform 1 0 1580 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2529
timestamp 1714281807
transform 1 0 1516 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2530
timestamp 1714281807
transform 1 0 1316 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2531
timestamp 1714281807
transform 1 0 1900 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2532
timestamp 1714281807
transform 1 0 1852 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2533
timestamp 1714281807
transform 1 0 1852 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2534
timestamp 1714281807
transform 1 0 1876 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2535
timestamp 1714281807
transform 1 0 1788 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2536
timestamp 1714281807
transform 1 0 1628 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2537
timestamp 1714281807
transform 1 0 1636 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2538
timestamp 1714281807
transform 1 0 1636 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2539
timestamp 1714281807
transform 1 0 1748 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2540
timestamp 1714281807
transform 1 0 1652 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2541
timestamp 1714281807
transform 1 0 1564 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2542
timestamp 1714281807
transform 1 0 1516 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2543
timestamp 1714281807
transform 1 0 1732 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2544
timestamp 1714281807
transform 1 0 1628 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2545
timestamp 1714281807
transform 1 0 668 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2546
timestamp 1714281807
transform 1 0 644 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_2547
timestamp 1714281807
transform 1 0 644 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2548
timestamp 1714281807
transform 1 0 324 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2549
timestamp 1714281807
transform 1 0 1204 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_2550
timestamp 1714281807
transform 1 0 1164 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2551
timestamp 1714281807
transform 1 0 1060 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2552
timestamp 1714281807
transform 1 0 1060 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_2553
timestamp 1714281807
transform 1 0 940 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2554
timestamp 1714281807
transform 1 0 836 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2555
timestamp 1714281807
transform 1 0 700 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2556
timestamp 1714281807
transform 1 0 652 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2557
timestamp 1714281807
transform 1 0 620 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_2558
timestamp 1714281807
transform 1 0 604 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2559
timestamp 1714281807
transform 1 0 516 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2560
timestamp 1714281807
transform 1 0 492 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2561
timestamp 1714281807
transform 1 0 476 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2562
timestamp 1714281807
transform 1 0 396 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2563
timestamp 1714281807
transform 1 0 420 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2564
timestamp 1714281807
transform 1 0 316 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2565
timestamp 1714281807
transform 1 0 308 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2566
timestamp 1714281807
transform 1 0 268 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2567
timestamp 1714281807
transform 1 0 268 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2568
timestamp 1714281807
transform 1 0 228 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2569
timestamp 1714281807
transform 1 0 204 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2570
timestamp 1714281807
transform 1 0 292 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2571
timestamp 1714281807
transform 1 0 236 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2572
timestamp 1714281807
transform 1 0 236 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2573
timestamp 1714281807
transform 1 0 692 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2574
timestamp 1714281807
transform 1 0 692 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2575
timestamp 1714281807
transform 1 0 340 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2576
timestamp 1714281807
transform 1 0 332 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2577
timestamp 1714281807
transform 1 0 316 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2578
timestamp 1714281807
transform 1 0 724 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2579
timestamp 1714281807
transform 1 0 684 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2580
timestamp 1714281807
transform 1 0 668 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2581
timestamp 1714281807
transform 1 0 780 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2582
timestamp 1714281807
transform 1 0 740 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2583
timestamp 1714281807
transform 1 0 844 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2584
timestamp 1714281807
transform 1 0 836 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2585
timestamp 1714281807
transform 1 0 756 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2586
timestamp 1714281807
transform 1 0 420 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2587
timestamp 1714281807
transform 1 0 220 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2588
timestamp 1714281807
transform 1 0 196 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2589
timestamp 1714281807
transform 1 0 740 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2590
timestamp 1714281807
transform 1 0 724 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2591
timestamp 1714281807
transform 1 0 740 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2592
timestamp 1714281807
transform 1 0 708 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2593
timestamp 1714281807
transform 1 0 572 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2594
timestamp 1714281807
transform 1 0 548 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2595
timestamp 1714281807
transform 1 0 492 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2596
timestamp 1714281807
transform 1 0 196 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2597
timestamp 1714281807
transform 1 0 644 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2598
timestamp 1714281807
transform 1 0 644 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2599
timestamp 1714281807
transform 1 0 692 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2600
timestamp 1714281807
transform 1 0 692 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2601
timestamp 1714281807
transform 1 0 884 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2602
timestamp 1714281807
transform 1 0 812 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2603
timestamp 1714281807
transform 1 0 804 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2604
timestamp 1714281807
transform 1 0 1060 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2605
timestamp 1714281807
transform 1 0 964 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2606
timestamp 1714281807
transform 1 0 1396 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2607
timestamp 1714281807
transform 1 0 1284 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2608
timestamp 1714281807
transform 1 0 748 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2609
timestamp 1714281807
transform 1 0 708 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2610
timestamp 1714281807
transform 1 0 708 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2611
timestamp 1714281807
transform 1 0 924 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_2612
timestamp 1714281807
transform 1 0 900 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2613
timestamp 1714281807
transform 1 0 980 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2614
timestamp 1714281807
transform 1 0 964 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_2615
timestamp 1714281807
transform 1 0 852 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2616
timestamp 1714281807
transform 1 0 844 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2617
timestamp 1714281807
transform 1 0 812 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2618
timestamp 1714281807
transform 1 0 1012 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2619
timestamp 1714281807
transform 1 0 996 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2620
timestamp 1714281807
transform 1 0 1028 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_2621
timestamp 1714281807
transform 1 0 1028 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2622
timestamp 1714281807
transform 1 0 1308 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2623
timestamp 1714281807
transform 1 0 1276 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2624
timestamp 1714281807
transform 1 0 1412 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2625
timestamp 1714281807
transform 1 0 1220 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2626
timestamp 1714281807
transform 1 0 1188 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_2627
timestamp 1714281807
transform 1 0 1308 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2628
timestamp 1714281807
transform 1 0 1260 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2629
timestamp 1714281807
transform 1 0 1404 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2630
timestamp 1714281807
transform 1 0 1228 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2631
timestamp 1714281807
transform 1 0 1932 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2632
timestamp 1714281807
transform 1 0 1868 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2633
timestamp 1714281807
transform 1 0 1860 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2634
timestamp 1714281807
transform 1 0 1844 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_2635
timestamp 1714281807
transform 1 0 1460 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2636
timestamp 1714281807
transform 1 0 1380 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2637
timestamp 1714281807
transform 1 0 2524 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2638
timestamp 1714281807
transform 1 0 2492 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2639
timestamp 1714281807
transform 1 0 2604 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2640
timestamp 1714281807
transform 1 0 2588 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2641
timestamp 1714281807
transform 1 0 2324 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2642
timestamp 1714281807
transform 1 0 2316 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2643
timestamp 1714281807
transform 1 0 2156 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2644
timestamp 1714281807
transform 1 0 2148 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2645
timestamp 1714281807
transform 1 0 2068 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2646
timestamp 1714281807
transform 1 0 2012 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2647
timestamp 1714281807
transform 1 0 1892 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2648
timestamp 1714281807
transform 1 0 1892 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2649
timestamp 1714281807
transform 1 0 1556 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2650
timestamp 1714281807
transform 1 0 1540 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2651
timestamp 1714281807
transform 1 0 1708 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2652
timestamp 1714281807
transform 1 0 1700 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2653
timestamp 1714281807
transform 1 0 1452 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2654
timestamp 1714281807
transform 1 0 1436 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2655
timestamp 1714281807
transform 1 0 1084 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2656
timestamp 1714281807
transform 1 0 988 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2657
timestamp 1714281807
transform 1 0 1132 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2658
timestamp 1714281807
transform 1 0 1108 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2659
timestamp 1714281807
transform 1 0 1300 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2660
timestamp 1714281807
transform 1 0 1300 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2661
timestamp 1714281807
transform 1 0 1132 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2662
timestamp 1714281807
transform 1 0 1028 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2663
timestamp 1714281807
transform 1 0 1116 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2664
timestamp 1714281807
transform 1 0 1020 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2665
timestamp 1714281807
transform 1 0 1308 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2666
timestamp 1714281807
transform 1 0 1228 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2667
timestamp 1714281807
transform 1 0 1876 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2668
timestamp 1714281807
transform 1 0 1876 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2669
timestamp 1714281807
transform 1 0 1636 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2670
timestamp 1714281807
transform 1 0 1636 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2671
timestamp 1714281807
transform 1 0 1900 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2672
timestamp 1714281807
transform 1 0 1884 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2673
timestamp 1714281807
transform 1 0 1580 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2674
timestamp 1714281807
transform 1 0 1572 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2675
timestamp 1714281807
transform 1 0 1588 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2676
timestamp 1714281807
transform 1 0 1572 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2677
timestamp 1714281807
transform 1 0 1836 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2678
timestamp 1714281807
transform 1 0 1796 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2679
timestamp 1714281807
transform 1 0 2460 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2680
timestamp 1714281807
transform 1 0 2420 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2681
timestamp 1714281807
transform 1 0 2460 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2682
timestamp 1714281807
transform 1 0 2452 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2683
timestamp 1714281807
transform 1 0 2436 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2684
timestamp 1714281807
transform 1 0 2396 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2685
timestamp 1714281807
transform 1 0 2940 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2686
timestamp 1714281807
transform 1 0 2868 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2687
timestamp 1714281807
transform 1 0 2804 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2688
timestamp 1714281807
transform 1 0 2804 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2689
timestamp 1714281807
transform 1 0 2908 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2690
timestamp 1714281807
transform 1 0 2900 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2691
timestamp 1714281807
transform 1 0 2316 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2692
timestamp 1714281807
transform 1 0 2308 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2693
timestamp 1714281807
transform 1 0 2156 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2694
timestamp 1714281807
transform 1 0 2092 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2695
timestamp 1714281807
transform 1 0 2444 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2696
timestamp 1714281807
transform 1 0 2436 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2697
timestamp 1714281807
transform 1 0 1900 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2698
timestamp 1714281807
transform 1 0 1868 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2699
timestamp 1714281807
transform 1 0 1788 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2700
timestamp 1714281807
transform 1 0 1756 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2701
timestamp 1714281807
transform 1 0 1988 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2702
timestamp 1714281807
transform 1 0 1980 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2703
timestamp 1714281807
transform 1 0 2796 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2704
timestamp 1714281807
transform 1 0 2796 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2705
timestamp 1714281807
transform 1 0 2532 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2706
timestamp 1714281807
transform 1 0 2532 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2707
timestamp 1714281807
transform 1 0 2916 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2708
timestamp 1714281807
transform 1 0 2852 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2709
timestamp 1714281807
transform 1 0 1324 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_2710
timestamp 1714281807
transform 1 0 1316 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2711
timestamp 1714281807
transform 1 0 1468 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_2712
timestamp 1714281807
transform 1 0 1436 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2713
timestamp 1714281807
transform 1 0 1404 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_2714
timestamp 1714281807
transform 1 0 1332 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2715
timestamp 1714281807
transform 1 0 2940 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2716
timestamp 1714281807
transform 1 0 2860 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2717
timestamp 1714281807
transform 1 0 2652 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2718
timestamp 1714281807
transform 1 0 2644 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2719
timestamp 1714281807
transform 1 0 2924 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2720
timestamp 1714281807
transform 1 0 2884 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2721
timestamp 1714281807
transform 1 0 2372 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_2722
timestamp 1714281807
transform 1 0 2292 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2723
timestamp 1714281807
transform 1 0 2172 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2724
timestamp 1714281807
transform 1 0 2172 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2725
timestamp 1714281807
transform 1 0 2340 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2726
timestamp 1714281807
transform 1 0 2260 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2727
timestamp 1714281807
transform 1 0 2940 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2728
timestamp 1714281807
transform 1 0 2868 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2729
timestamp 1714281807
transform 1 0 2772 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2730
timestamp 1714281807
transform 1 0 2772 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2731
timestamp 1714281807
transform 1 0 2940 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2732
timestamp 1714281807
transform 1 0 2868 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2733
timestamp 1714281807
transform 1 0 452 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2734
timestamp 1714281807
transform 1 0 372 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2735
timestamp 1714281807
transform 1 0 524 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2736
timestamp 1714281807
transform 1 0 484 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2737
timestamp 1714281807
transform 1 0 604 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2738
timestamp 1714281807
transform 1 0 596 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2739
timestamp 1714281807
transform 1 0 772 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2740
timestamp 1714281807
transform 1 0 692 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2741
timestamp 1714281807
transform 1 0 540 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2742
timestamp 1714281807
transform 1 0 396 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2743
timestamp 1714281807
transform 1 0 548 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2744
timestamp 1714281807
transform 1 0 396 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2745
timestamp 1714281807
transform 1 0 2444 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2746
timestamp 1714281807
transform 1 0 2444 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2747
timestamp 1714281807
transform 1 0 2468 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2748
timestamp 1714281807
transform 1 0 2364 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2749
timestamp 1714281807
transform 1 0 2380 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2750
timestamp 1714281807
transform 1 0 2316 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2751
timestamp 1714281807
transform 1 0 2428 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2752
timestamp 1714281807
transform 1 0 2428 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2753
timestamp 1714281807
transform 1 0 2508 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2754
timestamp 1714281807
transform 1 0 2508 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2755
timestamp 1714281807
transform 1 0 2340 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2756
timestamp 1714281807
transform 1 0 2324 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2757
timestamp 1714281807
transform 1 0 2044 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2758
timestamp 1714281807
transform 1 0 1980 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2759
timestamp 1714281807
transform 1 0 2172 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2760
timestamp 1714281807
transform 1 0 2164 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2761
timestamp 1714281807
transform 1 0 1852 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2762
timestamp 1714281807
transform 1 0 1844 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2763
timestamp 1714281807
transform 1 0 1780 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2764
timestamp 1714281807
transform 1 0 1780 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2765
timestamp 1714281807
transform 1 0 1988 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2766
timestamp 1714281807
transform 1 0 1948 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2767
timestamp 1714281807
transform 1 0 1884 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2768
timestamp 1714281807
transform 1 0 1860 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2769
timestamp 1714281807
transform 1 0 1436 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2770
timestamp 1714281807
transform 1 0 1316 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2771
timestamp 1714281807
transform 1 0 1700 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2772
timestamp 1714281807
transform 1 0 1644 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2773
timestamp 1714281807
transform 1 0 1444 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2774
timestamp 1714281807
transform 1 0 1308 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2775
timestamp 1714281807
transform 1 0 1452 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2776
timestamp 1714281807
transform 1 0 1452 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2777
timestamp 1714281807
transform 1 0 1572 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2778
timestamp 1714281807
transform 1 0 1492 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2779
timestamp 1714281807
transform 1 0 1524 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2780
timestamp 1714281807
transform 1 0 1508 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2781
timestamp 1714281807
transform 1 0 1468 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2782
timestamp 1714281807
transform 1 0 1372 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2783
timestamp 1714281807
transform 1 0 1412 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2784
timestamp 1714281807
transform 1 0 1300 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2785
timestamp 1714281807
transform 1 0 1556 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2786
timestamp 1714281807
transform 1 0 1476 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2787
timestamp 1714281807
transform 1 0 2020 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2788
timestamp 1714281807
transform 1 0 1940 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2789
timestamp 1714281807
transform 1 0 1988 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2790
timestamp 1714281807
transform 1 0 1988 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2791
timestamp 1714281807
transform 1 0 2028 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2792
timestamp 1714281807
transform 1 0 1948 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2793
timestamp 1714281807
transform 1 0 2164 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2794
timestamp 1714281807
transform 1 0 2076 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2795
timestamp 1714281807
transform 1 0 2108 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2796
timestamp 1714281807
transform 1 0 2020 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2797
timestamp 1714281807
transform 1 0 2004 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2798
timestamp 1714281807
transform 1 0 1964 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2799
timestamp 1714281807
transform 1 0 2724 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2800
timestamp 1714281807
transform 1 0 2724 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2801
timestamp 1714281807
transform 1 0 2628 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2802
timestamp 1714281807
transform 1 0 2628 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2803
timestamp 1714281807
transform 1 0 2492 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2804
timestamp 1714281807
transform 1 0 2484 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2805
timestamp 1714281807
transform 1 0 2644 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2806
timestamp 1714281807
transform 1 0 2644 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2807
timestamp 1714281807
transform 1 0 2716 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2808
timestamp 1714281807
transform 1 0 2676 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2809
timestamp 1714281807
transform 1 0 2524 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2810
timestamp 1714281807
transform 1 0 2524 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2811
timestamp 1714281807
transform 1 0 1988 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2812
timestamp 1714281807
transform 1 0 1908 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2813
timestamp 1714281807
transform 1 0 1900 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2814
timestamp 1714281807
transform 1 0 1892 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2815
timestamp 1714281807
transform 1 0 1812 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2816
timestamp 1714281807
transform 1 0 1804 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2817
timestamp 1714281807
transform 1 0 2356 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2818
timestamp 1714281807
transform 1 0 2348 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2819
timestamp 1714281807
transform 1 0 2236 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2820
timestamp 1714281807
transform 1 0 2228 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2821
timestamp 1714281807
transform 1 0 2148 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2822
timestamp 1714281807
transform 1 0 2132 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2823
timestamp 1714281807
transform 1 0 2764 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2824
timestamp 1714281807
transform 1 0 2700 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2825
timestamp 1714281807
transform 1 0 2796 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2826
timestamp 1714281807
transform 1 0 2796 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2827
timestamp 1714281807
transform 1 0 2700 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2828
timestamp 1714281807
transform 1 0 2700 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2829
timestamp 1714281807
transform 1 0 2428 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2830
timestamp 1714281807
transform 1 0 2388 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2831
timestamp 1714281807
transform 1 0 2172 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2832
timestamp 1714281807
transform 1 0 2172 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2833
timestamp 1714281807
transform 1 0 2236 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2834
timestamp 1714281807
transform 1 0 2188 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2835
timestamp 1714281807
transform 1 0 604 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2836
timestamp 1714281807
transform 1 0 596 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2837
timestamp 1714281807
transform 1 0 468 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2838
timestamp 1714281807
transform 1 0 372 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2839
timestamp 1714281807
transform 1 0 420 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2840
timestamp 1714281807
transform 1 0 420 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2841
timestamp 1714281807
transform 1 0 324 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2842
timestamp 1714281807
transform 1 0 284 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2843
timestamp 1714281807
transform 1 0 300 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2844
timestamp 1714281807
transform 1 0 156 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2845
timestamp 1714281807
transform 1 0 340 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2846
timestamp 1714281807
transform 1 0 188 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2847
timestamp 1714281807
transform 1 0 420 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2848
timestamp 1714281807
transform 1 0 324 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2849
timestamp 1714281807
transform 1 0 580 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2850
timestamp 1714281807
transform 1 0 556 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2851
timestamp 1714281807
transform 1 0 884 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2852
timestamp 1714281807
transform 1 0 828 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2853
timestamp 1714281807
transform 1 0 1324 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2854
timestamp 1714281807
transform 1 0 1284 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2855
timestamp 1714281807
transform 1 0 756 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2856
timestamp 1714281807
transform 1 0 748 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2857
timestamp 1714281807
transform 1 0 860 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2858
timestamp 1714281807
transform 1 0 860 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2859
timestamp 1714281807
transform 1 0 1332 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2860
timestamp 1714281807
transform 1 0 1332 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2861
timestamp 1714281807
transform 1 0 1164 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2862
timestamp 1714281807
transform 1 0 1148 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2863
timestamp 1714281807
transform 1 0 1196 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2864
timestamp 1714281807
transform 1 0 1108 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2865
timestamp 1714281807
transform 1 0 1164 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2866
timestamp 1714281807
transform 1 0 1076 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2867
timestamp 1714281807
transform 1 0 2756 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2868
timestamp 1714281807
transform 1 0 2676 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2869
timestamp 1714281807
transform 1 0 2748 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2870
timestamp 1714281807
transform 1 0 2660 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2871
timestamp 1714281807
transform 1 0 2732 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2872
timestamp 1714281807
transform 1 0 2644 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2873
timestamp 1714281807
transform 1 0 860 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2874
timestamp 1714281807
transform 1 0 820 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2875
timestamp 1714281807
transform 1 0 604 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2876
timestamp 1714281807
transform 1 0 556 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2877
timestamp 1714281807
transform 1 0 460 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2878
timestamp 1714281807
transform 1 0 412 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2879
timestamp 1714281807
transform 1 0 396 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2880
timestamp 1714281807
transform 1 0 396 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2881
timestamp 1714281807
transform 1 0 580 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2882
timestamp 1714281807
transform 1 0 580 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2883
timestamp 1714281807
transform 1 0 692 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2884
timestamp 1714281807
transform 1 0 692 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2885
timestamp 1714281807
transform 1 0 476 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2886
timestamp 1714281807
transform 1 0 476 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2887
timestamp 1714281807
transform 1 0 788 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2888
timestamp 1714281807
transform 1 0 788 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2889
timestamp 1714281807
transform 1 0 876 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2890
timestamp 1714281807
transform 1 0 876 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2891
timestamp 1714281807
transform 1 0 884 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2892
timestamp 1714281807
transform 1 0 860 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2893
timestamp 1714281807
transform 1 0 788 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2894
timestamp 1714281807
transform 1 0 652 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2895
timestamp 1714281807
transform 1 0 636 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2896
timestamp 1714281807
transform 1 0 812 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2897
timestamp 1714281807
transform 1 0 796 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_2898
timestamp 1714281807
transform 1 0 764 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_2899
timestamp 1714281807
transform 1 0 764 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2900
timestamp 1714281807
transform 1 0 636 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2901
timestamp 1714281807
transform 1 0 548 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2902
timestamp 1714281807
transform 1 0 356 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2903
timestamp 1714281807
transform 1 0 356 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2904
timestamp 1714281807
transform 1 0 428 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2905
timestamp 1714281807
transform 1 0 420 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2906
timestamp 1714281807
transform 1 0 404 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2907
timestamp 1714281807
transform 1 0 684 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2908
timestamp 1714281807
transform 1 0 660 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2909
timestamp 1714281807
transform 1 0 636 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2910
timestamp 1714281807
transform 1 0 636 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2911
timestamp 1714281807
transform 1 0 604 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2912
timestamp 1714281807
transform 1 0 604 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2913
timestamp 1714281807
transform 1 0 780 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2914
timestamp 1714281807
transform 1 0 692 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2915
timestamp 1714281807
transform 1 0 676 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2916
timestamp 1714281807
transform 1 0 588 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2917
timestamp 1714281807
transform 1 0 564 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2918
timestamp 1714281807
transform 1 0 492 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2919
timestamp 1714281807
transform 1 0 540 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2920
timestamp 1714281807
transform 1 0 540 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2921
timestamp 1714281807
transform 1 0 676 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2922
timestamp 1714281807
transform 1 0 572 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2923
timestamp 1714281807
transform 1 0 572 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2924
timestamp 1714281807
transform 1 0 548 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_2925
timestamp 1714281807
transform 1 0 316 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2926
timestamp 1714281807
transform 1 0 284 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2927
timestamp 1714281807
transform 1 0 620 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_2928
timestamp 1714281807
transform 1 0 444 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_2929
timestamp 1714281807
transform 1 0 428 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2930
timestamp 1714281807
transform 1 0 412 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2931
timestamp 1714281807
transform 1 0 844 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2932
timestamp 1714281807
transform 1 0 844 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2933
timestamp 1714281807
transform 1 0 652 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2934
timestamp 1714281807
transform 1 0 436 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2935
timestamp 1714281807
transform 1 0 708 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2936
timestamp 1714281807
transform 1 0 684 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2937
timestamp 1714281807
transform 1 0 780 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2938
timestamp 1714281807
transform 1 0 692 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2939
timestamp 1714281807
transform 1 0 708 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2940
timestamp 1714281807
transform 1 0 676 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2941
timestamp 1714281807
transform 1 0 508 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2942
timestamp 1714281807
transform 1 0 356 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2943
timestamp 1714281807
transform 1 0 524 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2944
timestamp 1714281807
transform 1 0 476 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2945
timestamp 1714281807
transform 1 0 500 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2946
timestamp 1714281807
transform 1 0 484 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2947
timestamp 1714281807
transform 1 0 500 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2948
timestamp 1714281807
transform 1 0 500 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2949
timestamp 1714281807
transform 1 0 444 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_2950
timestamp 1714281807
transform 1 0 412 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2951
timestamp 1714281807
transform 1 0 580 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2952
timestamp 1714281807
transform 1 0 548 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2953
timestamp 1714281807
transform 1 0 788 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2954
timestamp 1714281807
transform 1 0 508 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2955
timestamp 1714281807
transform 1 0 516 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2956
timestamp 1714281807
transform 1 0 508 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2957
timestamp 1714281807
transform 1 0 500 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2958
timestamp 1714281807
transform 1 0 516 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2959
timestamp 1714281807
transform 1 0 396 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2960
timestamp 1714281807
transform 1 0 524 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2961
timestamp 1714281807
transform 1 0 460 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2962
timestamp 1714281807
transform 1 0 428 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2963
timestamp 1714281807
transform 1 0 428 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_2964
timestamp 1714281807
transform 1 0 372 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2965
timestamp 1714281807
transform 1 0 308 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2966
timestamp 1714281807
transform 1 0 868 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_2967
timestamp 1714281807
transform 1 0 868 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2968
timestamp 1714281807
transform 1 0 2052 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_2969
timestamp 1714281807
transform 1 0 1996 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_2970
timestamp 1714281807
transform 1 0 1860 0 1 1585
box -2 -2 2 2
use M2_M1  M2_M1_2971
timestamp 1714281807
transform 1 0 1812 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_2972
timestamp 1714281807
transform 1 0 1756 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_2973
timestamp 1714281807
transform 1 0 1756 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_2974
timestamp 1714281807
transform 1 0 1716 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_2975
timestamp 1714281807
transform 1 0 1668 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_2976
timestamp 1714281807
transform 1 0 1668 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_2977
timestamp 1714281807
transform 1 0 1668 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_2978
timestamp 1714281807
transform 1 0 1580 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_2979
timestamp 1714281807
transform 1 0 1540 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_2980
timestamp 1714281807
transform 1 0 1436 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_2981
timestamp 1714281807
transform 1 0 1076 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_2982
timestamp 1714281807
transform 1 0 1036 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2983
timestamp 1714281807
transform 1 0 1036 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_2984
timestamp 1714281807
transform 1 0 948 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2985
timestamp 1714281807
transform 1 0 756 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2986
timestamp 1714281807
transform 1 0 748 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2987
timestamp 1714281807
transform 1 0 780 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_2988
timestamp 1714281807
transform 1 0 548 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2989
timestamp 1714281807
transform 1 0 524 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_2990
timestamp 1714281807
transform 1 0 492 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2991
timestamp 1714281807
transform 1 0 828 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2992
timestamp 1714281807
transform 1 0 740 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2993
timestamp 1714281807
transform 1 0 756 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_2994
timestamp 1714281807
transform 1 0 724 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_2995
timestamp 1714281807
transform 1 0 892 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_2996
timestamp 1714281807
transform 1 0 668 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_2997
timestamp 1714281807
transform 1 0 892 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2998
timestamp 1714281807
transform 1 0 836 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_2999
timestamp 1714281807
transform 1 0 756 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3000
timestamp 1714281807
transform 1 0 732 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_3001
timestamp 1714281807
transform 1 0 500 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_3002
timestamp 1714281807
transform 1 0 260 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3003
timestamp 1714281807
transform 1 0 812 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3004
timestamp 1714281807
transform 1 0 796 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3005
timestamp 1714281807
transform 1 0 564 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3006
timestamp 1714281807
transform 1 0 564 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3007
timestamp 1714281807
transform 1 0 644 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_3008
timestamp 1714281807
transform 1 0 516 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_3009
timestamp 1714281807
transform 1 0 404 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_3010
timestamp 1714281807
transform 1 0 708 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3011
timestamp 1714281807
transform 1 0 708 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3012
timestamp 1714281807
transform 1 0 612 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3013
timestamp 1714281807
transform 1 0 460 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3014
timestamp 1714281807
transform 1 0 2268 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3015
timestamp 1714281807
transform 1 0 2092 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3016
timestamp 1714281807
transform 1 0 2212 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3017
timestamp 1714281807
transform 1 0 2964 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3018
timestamp 1714281807
transform 1 0 2956 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3019
timestamp 1714281807
transform 1 0 3012 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3020
timestamp 1714281807
transform 1 0 2460 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3021
timestamp 1714281807
transform 1 0 2324 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3022
timestamp 1714281807
transform 1 0 2164 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3023
timestamp 1714281807
transform 1 0 2068 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3024
timestamp 1714281807
transform 1 0 2100 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3025
timestamp 1714281807
transform 1 0 1836 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3026
timestamp 1714281807
transform 1 0 2964 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3027
timestamp 1714281807
transform 1 0 2908 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3028
timestamp 1714281807
transform 1 0 2564 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3029
timestamp 1714281807
transform 1 0 1700 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3030
timestamp 1714281807
transform 1 0 1740 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3031
timestamp 1714281807
transform 1 0 1708 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3032
timestamp 1714281807
transform 1 0 3012 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3033
timestamp 1714281807
transform 1 0 2964 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3034
timestamp 1714281807
transform 1 0 2636 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3035
timestamp 1714281807
transform 1 0 2404 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3036
timestamp 1714281807
transform 1 0 2676 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3037
timestamp 1714281807
transform 1 0 2220 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3038
timestamp 1714281807
transform 1 0 2940 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3039
timestamp 1714281807
transform 1 0 2948 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3040
timestamp 1714281807
transform 1 0 2988 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3041
timestamp 1714281807
transform 1 0 2668 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3042
timestamp 1714281807
transform 1 0 2660 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3043
timestamp 1714281807
transform 1 0 2436 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3044
timestamp 1714281807
transform 1 0 2308 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3045
timestamp 1714281807
transform 1 0 2292 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3046
timestamp 1714281807
transform 1 0 1932 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3047
timestamp 1714281807
transform 1 0 1652 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3048
timestamp 1714281807
transform 1 0 2164 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3049
timestamp 1714281807
transform 1 0 2108 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3050
timestamp 1714281807
transform 1 0 1628 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3051
timestamp 1714281807
transform 1 0 1748 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3052
timestamp 1714281807
transform 1 0 1604 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3053
timestamp 1714281807
transform 1 0 1620 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3054
timestamp 1714281807
transform 1 0 1556 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3055
timestamp 1714281807
transform 1 0 1604 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3056
timestamp 1714281807
transform 1 0 2132 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3057
timestamp 1714281807
transform 1 0 2228 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3058
timestamp 1714281807
transform 1 0 2188 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3059
timestamp 1714281807
transform 1 0 2276 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3060
timestamp 1714281807
transform 1 0 2324 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3061
timestamp 1714281807
transform 1 0 1956 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3062
timestamp 1714281807
transform 1 0 2596 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3063
timestamp 1714281807
transform 1 0 2580 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3064
timestamp 1714281807
transform 1 0 2588 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3065
timestamp 1714281807
transform 1 0 2636 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3066
timestamp 1714281807
transform 1 0 2588 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3067
timestamp 1714281807
transform 1 0 2676 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3068
timestamp 1714281807
transform 1 0 2556 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3069
timestamp 1714281807
transform 1 0 2388 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3070
timestamp 1714281807
transform 1 0 2220 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3071
timestamp 1714281807
transform 1 0 2068 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3072
timestamp 1714281807
transform 1 0 1972 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3073
timestamp 1714281807
transform 1 0 1764 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3074
timestamp 1714281807
transform 1 0 2868 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3075
timestamp 1714281807
transform 1 0 2772 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3076
timestamp 1714281807
transform 1 0 2660 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3077
timestamp 1714281807
transform 1 0 1692 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3078
timestamp 1714281807
transform 1 0 1748 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3079
timestamp 1714281807
transform 1 0 1660 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3080
timestamp 1714281807
transform 1 0 3012 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3081
timestamp 1714281807
transform 1 0 2828 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3082
timestamp 1714281807
transform 1 0 2676 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3083
timestamp 1714281807
transform 1 0 2580 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3084
timestamp 1714281807
transform 1 0 2572 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3085
timestamp 1714281807
transform 1 0 2740 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3086
timestamp 1714281807
transform 1 0 2996 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3087
timestamp 1714281807
transform 1 0 2996 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3088
timestamp 1714281807
transform 1 0 2844 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3089
timestamp 1714281807
transform 1 0 2564 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3090
timestamp 1714281807
transform 1 0 2708 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3091
timestamp 1714281807
transform 1 0 2388 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3092
timestamp 1714281807
transform 1 0 2220 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3093
timestamp 1714281807
transform 1 0 1980 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3094
timestamp 1714281807
transform 1 0 1828 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3095
timestamp 1714281807
transform 1 0 1508 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3096
timestamp 1714281807
transform 1 0 1668 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3097
timestamp 1714281807
transform 1 0 1332 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3098
timestamp 1714281807
transform 1 0 1020 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3099
timestamp 1714281807
transform 1 0 1036 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3100
timestamp 1714281807
transform 1 0 1148 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3101
timestamp 1714281807
transform 1 0 1004 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3102
timestamp 1714281807
transform 1 0 996 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3103
timestamp 1714281807
transform 1 0 1156 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3104
timestamp 1714281807
transform 1 0 1836 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3105
timestamp 1714281807
transform 1 0 1716 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3106
timestamp 1714281807
transform 1 0 1852 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3107
timestamp 1714281807
transform 1 0 1700 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3108
timestamp 1714281807
transform 1 0 1668 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3109
timestamp 1714281807
transform 1 0 1804 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3110
timestamp 1714281807
transform 1 0 324 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3111
timestamp 1714281807
transform 1 0 356 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3112
timestamp 1714281807
transform 1 0 292 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3113
timestamp 1714281807
transform 1 0 244 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3114
timestamp 1714281807
transform 1 0 332 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3115
timestamp 1714281807
transform 1 0 308 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3116
timestamp 1714281807
transform 1 0 220 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3117
timestamp 1714281807
transform 1 0 180 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3118
timestamp 1714281807
transform 1 0 796 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3119
timestamp 1714281807
transform 1 0 1508 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3120
timestamp 1714281807
transform 1 0 804 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3121
timestamp 1714281807
transform 1 0 828 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3122
timestamp 1714281807
transform 1 0 1484 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3123
timestamp 1714281807
transform 1 0 1548 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3124
timestamp 1714281807
transform 1 0 1476 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3125
timestamp 1714281807
transform 1 0 1468 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3126
timestamp 1714281807
transform 1 0 940 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3127
timestamp 1714281807
transform 1 0 908 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3128
timestamp 1714281807
transform 1 0 916 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3129
timestamp 1714281807
transform 1 0 876 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_3130
timestamp 1714281807
transform 1 0 828 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_3131
timestamp 1714281807
transform 1 0 804 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_3132
timestamp 1714281807
transform 1 0 820 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3133
timestamp 1714281807
transform 1 0 820 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3134
timestamp 1714281807
transform 1 0 732 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3135
timestamp 1714281807
transform 1 0 676 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3136
timestamp 1714281807
transform 1 0 620 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3137
timestamp 1714281807
transform 1 0 532 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3138
timestamp 1714281807
transform 1 0 436 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3139
timestamp 1714281807
transform 1 0 724 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3140
timestamp 1714281807
transform 1 0 700 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3141
timestamp 1714281807
transform 1 0 692 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_3142
timestamp 1714281807
transform 1 0 628 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3143
timestamp 1714281807
transform 1 0 628 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3144
timestamp 1714281807
transform 1 0 436 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3145
timestamp 1714281807
transform 1 0 420 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_3146
timestamp 1714281807
transform 1 0 1052 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3147
timestamp 1714281807
transform 1 0 1044 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3148
timestamp 1714281807
transform 1 0 1020 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3149
timestamp 1714281807
transform 1 0 988 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3150
timestamp 1714281807
transform 1 0 980 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3151
timestamp 1714281807
transform 1 0 972 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_3152
timestamp 1714281807
transform 1 0 916 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3153
timestamp 1714281807
transform 1 0 900 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3154
timestamp 1714281807
transform 1 0 876 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3155
timestamp 1714281807
transform 1 0 876 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3156
timestamp 1714281807
transform 1 0 1180 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_3157
timestamp 1714281807
transform 1 0 1164 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3158
timestamp 1714281807
transform 1 0 1084 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3159
timestamp 1714281807
transform 1 0 1060 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_3160
timestamp 1714281807
transform 1 0 1196 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3161
timestamp 1714281807
transform 1 0 1132 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3162
timestamp 1714281807
transform 1 0 1132 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_3163
timestamp 1714281807
transform 1 0 1068 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_3164
timestamp 1714281807
transform 1 0 1068 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_3165
timestamp 1714281807
transform 1 0 596 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3166
timestamp 1714281807
transform 1 0 580 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_3167
timestamp 1714281807
transform 1 0 580 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3168
timestamp 1714281807
transform 1 0 428 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3169
timestamp 1714281807
transform 1 0 572 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3170
timestamp 1714281807
transform 1 0 564 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3171
timestamp 1714281807
transform 1 0 524 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3172
timestamp 1714281807
transform 1 0 516 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_3173
timestamp 1714281807
transform 1 0 500 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_3174
timestamp 1714281807
transform 1 0 444 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_3175
timestamp 1714281807
transform 1 0 692 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3176
timestamp 1714281807
transform 1 0 660 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_3177
timestamp 1714281807
transform 1 0 620 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3178
timestamp 1714281807
transform 1 0 612 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3179
timestamp 1714281807
transform 1 0 572 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3180
timestamp 1714281807
transform 1 0 700 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_3181
timestamp 1714281807
transform 1 0 660 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3182
timestamp 1714281807
transform 1 0 596 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3183
timestamp 1714281807
transform 1 0 1652 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3184
timestamp 1714281807
transform 1 0 1628 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3185
timestamp 1714281807
transform 1 0 1588 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3186
timestamp 1714281807
transform 1 0 1388 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3187
timestamp 1714281807
transform 1 0 1756 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3188
timestamp 1714281807
transform 1 0 1732 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3189
timestamp 1714281807
transform 1 0 1620 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3190
timestamp 1714281807
transform 1 0 1412 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3191
timestamp 1714281807
transform 1 0 1996 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3192
timestamp 1714281807
transform 1 0 1932 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3193
timestamp 1714281807
transform 1 0 1900 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3194
timestamp 1714281807
transform 1 0 1884 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3195
timestamp 1714281807
transform 1 0 1756 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3196
timestamp 1714281807
transform 1 0 1708 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3197
timestamp 1714281807
transform 1 0 1644 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3198
timestamp 1714281807
transform 1 0 1492 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_3199
timestamp 1714281807
transform 1 0 1292 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3200
timestamp 1714281807
transform 1 0 1628 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3201
timestamp 1714281807
transform 1 0 1572 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3202
timestamp 1714281807
transform 1 0 1564 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3203
timestamp 1714281807
transform 1 0 1484 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3204
timestamp 1714281807
transform 1 0 1276 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_3205
timestamp 1714281807
transform 1 0 892 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3206
timestamp 1714281807
transform 1 0 860 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3207
timestamp 1714281807
transform 1 0 764 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3208
timestamp 1714281807
transform 1 0 764 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3209
timestamp 1714281807
transform 1 0 628 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3210
timestamp 1714281807
transform 1 0 556 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3211
timestamp 1714281807
transform 1 0 372 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3212
timestamp 1714281807
transform 1 0 332 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3213
timestamp 1714281807
transform 1 0 780 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3214
timestamp 1714281807
transform 1 0 700 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3215
timestamp 1714281807
transform 1 0 684 0 1 105
box -2 -2 2 2
use M2_M1  M2_M1_3216
timestamp 1714281807
transform 1 0 628 0 1 105
box -2 -2 2 2
use M2_M1  M2_M1_3217
timestamp 1714281807
transform 1 0 548 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3218
timestamp 1714281807
transform 1 0 364 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3219
timestamp 1714281807
transform 1 0 348 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3220
timestamp 1714281807
transform 1 0 276 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3221
timestamp 1714281807
transform 1 0 220 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_3222
timestamp 1714281807
transform 1 0 620 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3223
timestamp 1714281807
transform 1 0 620 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_3224
timestamp 1714281807
transform 1 0 620 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3225
timestamp 1714281807
transform 1 0 588 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3226
timestamp 1714281807
transform 1 0 332 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3227
timestamp 1714281807
transform 1 0 324 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3228
timestamp 1714281807
transform 1 0 324 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_3229
timestamp 1714281807
transform 1 0 812 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3230
timestamp 1714281807
transform 1 0 812 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3231
timestamp 1714281807
transform 1 0 772 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3232
timestamp 1714281807
transform 1 0 660 0 1 185
box -2 -2 2 2
use M2_M1  M2_M1_3233
timestamp 1714281807
transform 1 0 380 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3234
timestamp 1714281807
transform 1 0 348 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3235
timestamp 1714281807
transform 1 0 260 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_3236
timestamp 1714281807
transform 1 0 260 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_3237
timestamp 1714281807
transform 1 0 1012 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3238
timestamp 1714281807
transform 1 0 844 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3239
timestamp 1714281807
transform 1 0 756 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3240
timestamp 1714281807
transform 1 0 892 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_3241
timestamp 1714281807
transform 1 0 812 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3242
timestamp 1714281807
transform 1 0 796 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3243
timestamp 1714281807
transform 1 0 780 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3244
timestamp 1714281807
transform 1 0 708 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3245
timestamp 1714281807
transform 1 0 876 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3246
timestamp 1714281807
transform 1 0 860 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3247
timestamp 1714281807
transform 1 0 340 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3248
timestamp 1714281807
transform 1 0 324 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3249
timestamp 1714281807
transform 1 0 300 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3250
timestamp 1714281807
transform 1 0 972 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_3251
timestamp 1714281807
transform 1 0 948 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_3252
timestamp 1714281807
transform 1 0 716 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3253
timestamp 1714281807
transform 1 0 508 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3254
timestamp 1714281807
transform 1 0 452 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3255
timestamp 1714281807
transform 1 0 420 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3256
timestamp 1714281807
transform 1 0 2036 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3257
timestamp 1714281807
transform 1 0 1708 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3258
timestamp 1714281807
transform 1 0 1476 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3259
timestamp 1714281807
transform 1 0 1004 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3260
timestamp 1714281807
transform 1 0 2916 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3261
timestamp 1714281807
transform 1 0 2916 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3262
timestamp 1714281807
transform 1 0 2916 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3263
timestamp 1714281807
transform 1 0 2916 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3264
timestamp 1714281807
transform 1 0 2900 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3265
timestamp 1714281807
transform 1 0 2892 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3266
timestamp 1714281807
transform 1 0 2868 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3267
timestamp 1714281807
transform 1 0 2780 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3268
timestamp 1714281807
transform 1 0 2772 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3269
timestamp 1714281807
transform 1 0 2764 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3270
timestamp 1714281807
transform 1 0 2724 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3271
timestamp 1714281807
transform 1 0 2692 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3272
timestamp 1714281807
transform 1 0 2676 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3273
timestamp 1714281807
transform 1 0 2676 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3274
timestamp 1714281807
transform 1 0 2652 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3275
timestamp 1714281807
transform 1 0 2628 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3276
timestamp 1714281807
transform 1 0 2612 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3277
timestamp 1714281807
transform 1 0 2612 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3278
timestamp 1714281807
transform 1 0 2596 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3279
timestamp 1714281807
transform 1 0 2596 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3280
timestamp 1714281807
transform 1 0 2580 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3281
timestamp 1714281807
transform 1 0 2540 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3282
timestamp 1714281807
transform 1 0 2500 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3283
timestamp 1714281807
transform 1 0 2492 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3284
timestamp 1714281807
transform 1 0 2460 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3285
timestamp 1714281807
transform 1 0 2444 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3286
timestamp 1714281807
transform 1 0 2444 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3287
timestamp 1714281807
transform 1 0 2436 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3288
timestamp 1714281807
transform 1 0 2420 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_3289
timestamp 1714281807
transform 1 0 2404 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3290
timestamp 1714281807
transform 1 0 2396 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3291
timestamp 1714281807
transform 1 0 2388 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3292
timestamp 1714281807
transform 1 0 2388 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3293
timestamp 1714281807
transform 1 0 2356 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3294
timestamp 1714281807
transform 1 0 2348 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3295
timestamp 1714281807
transform 1 0 2316 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3296
timestamp 1714281807
transform 1 0 2308 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3297
timestamp 1714281807
transform 1 0 2276 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3298
timestamp 1714281807
transform 1 0 2268 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3299
timestamp 1714281807
transform 1 0 2260 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3300
timestamp 1714281807
transform 1 0 2260 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3301
timestamp 1714281807
transform 1 0 2212 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3302
timestamp 1714281807
transform 1 0 2204 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3303
timestamp 1714281807
transform 1 0 2180 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3304
timestamp 1714281807
transform 1 0 2148 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3305
timestamp 1714281807
transform 1 0 2132 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3306
timestamp 1714281807
transform 1 0 2132 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3307
timestamp 1714281807
transform 1 0 2124 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3308
timestamp 1714281807
transform 1 0 2124 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3309
timestamp 1714281807
transform 1 0 2084 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3310
timestamp 1714281807
transform 1 0 2028 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3311
timestamp 1714281807
transform 1 0 1972 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3312
timestamp 1714281807
transform 1 0 1964 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3313
timestamp 1714281807
transform 1 0 1948 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3314
timestamp 1714281807
transform 1 0 1932 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3315
timestamp 1714281807
transform 1 0 1932 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3316
timestamp 1714281807
transform 1 0 1916 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3317
timestamp 1714281807
transform 1 0 1900 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3318
timestamp 1714281807
transform 1 0 1900 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3319
timestamp 1714281807
transform 1 0 1892 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3320
timestamp 1714281807
transform 1 0 1876 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3321
timestamp 1714281807
transform 1 0 1860 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3322
timestamp 1714281807
transform 1 0 1852 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3323
timestamp 1714281807
transform 1 0 1852 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3324
timestamp 1714281807
transform 1 0 1844 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3325
timestamp 1714281807
transform 1 0 1820 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3326
timestamp 1714281807
transform 1 0 1812 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3327
timestamp 1714281807
transform 1 0 1812 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3328
timestamp 1714281807
transform 1 0 1812 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3329
timestamp 1714281807
transform 1 0 1756 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3330
timestamp 1714281807
transform 1 0 1740 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3331
timestamp 1714281807
transform 1 0 1708 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3332
timestamp 1714281807
transform 1 0 1652 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3333
timestamp 1714281807
transform 1 0 1596 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3334
timestamp 1714281807
transform 1 0 1588 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3335
timestamp 1714281807
transform 1 0 1532 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3336
timestamp 1714281807
transform 1 0 1524 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3337
timestamp 1714281807
transform 1 0 1524 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3338
timestamp 1714281807
transform 1 0 1484 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3339
timestamp 1714281807
transform 1 0 1444 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3340
timestamp 1714281807
transform 1 0 1428 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3341
timestamp 1714281807
transform 1 0 1404 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3342
timestamp 1714281807
transform 1 0 1388 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3343
timestamp 1714281807
transform 1 0 1388 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3344
timestamp 1714281807
transform 1 0 1332 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3345
timestamp 1714281807
transform 1 0 1324 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3346
timestamp 1714281807
transform 1 0 1308 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3347
timestamp 1714281807
transform 1 0 1300 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3348
timestamp 1714281807
transform 1 0 1284 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3349
timestamp 1714281807
transform 1 0 1284 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3350
timestamp 1714281807
transform 1 0 1268 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3351
timestamp 1714281807
transform 1 0 1268 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3352
timestamp 1714281807
transform 1 0 1260 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3353
timestamp 1714281807
transform 1 0 1252 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3354
timestamp 1714281807
transform 1 0 1252 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3355
timestamp 1714281807
transform 1 0 1228 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3356
timestamp 1714281807
transform 1 0 1172 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3357
timestamp 1714281807
transform 1 0 1100 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3358
timestamp 1714281807
transform 1 0 1068 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3359
timestamp 1714281807
transform 1 0 1068 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3360
timestamp 1714281807
transform 1 0 1060 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3361
timestamp 1714281807
transform 1 0 1028 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3362
timestamp 1714281807
transform 1 0 1020 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3363
timestamp 1714281807
transform 1 0 980 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3364
timestamp 1714281807
transform 1 0 972 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3365
timestamp 1714281807
transform 1 0 972 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3366
timestamp 1714281807
transform 1 0 964 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3367
timestamp 1714281807
transform 1 0 948 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3368
timestamp 1714281807
transform 1 0 852 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3369
timestamp 1714281807
transform 1 0 836 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3370
timestamp 1714281807
transform 1 0 828 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3371
timestamp 1714281807
transform 1 0 796 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3372
timestamp 1714281807
transform 1 0 772 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3373
timestamp 1714281807
transform 1 0 756 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3374
timestamp 1714281807
transform 1 0 748 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3375
timestamp 1714281807
transform 1 0 700 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3376
timestamp 1714281807
transform 1 0 700 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3377
timestamp 1714281807
transform 1 0 692 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3378
timestamp 1714281807
transform 1 0 604 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3379
timestamp 1714281807
transform 1 0 572 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3380
timestamp 1714281807
transform 1 0 564 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_3381
timestamp 1714281807
transform 1 0 556 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3382
timestamp 1714281807
transform 1 0 556 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3383
timestamp 1714281807
transform 1 0 548 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3384
timestamp 1714281807
transform 1 0 508 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3385
timestamp 1714281807
transform 1 0 444 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3386
timestamp 1714281807
transform 1 0 436 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3387
timestamp 1714281807
transform 1 0 388 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3388
timestamp 1714281807
transform 1 0 372 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3389
timestamp 1714281807
transform 1 0 372 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3390
timestamp 1714281807
transform 1 0 372 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3391
timestamp 1714281807
transform 1 0 364 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3392
timestamp 1714281807
transform 1 0 332 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3393
timestamp 1714281807
transform 1 0 332 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3394
timestamp 1714281807
transform 1 0 324 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3395
timestamp 1714281807
transform 1 0 324 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3396
timestamp 1714281807
transform 1 0 308 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3397
timestamp 1714281807
transform 1 0 300 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3398
timestamp 1714281807
transform 1 0 276 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3399
timestamp 1714281807
transform 1 0 260 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3400
timestamp 1714281807
transform 1 0 196 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3401
timestamp 1714281807
transform 1 0 188 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_3402
timestamp 1714281807
transform 1 0 164 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3403
timestamp 1714281807
transform 1 0 140 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3404
timestamp 1714281807
transform 1 0 132 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3405
timestamp 1714281807
transform 1 0 108 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3406
timestamp 1714281807
transform 1 0 108 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_0
timestamp 1714281807
transform 1 0 1148 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_1
timestamp 1714281807
transform 1 0 948 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2
timestamp 1714281807
transform 1 0 860 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3
timestamp 1714281807
transform 1 0 836 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_4
timestamp 1714281807
transform 1 0 732 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_5
timestamp 1714281807
transform 1 0 628 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_6
timestamp 1714281807
transform 1 0 508 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_7
timestamp 1714281807
transform 1 0 604 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_8
timestamp 1714281807
transform 1 0 532 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_9
timestamp 1714281807
transform 1 0 780 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_10
timestamp 1714281807
transform 1 0 740 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_11
timestamp 1714281807
transform 1 0 932 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_12
timestamp 1714281807
transform 1 0 900 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_13
timestamp 1714281807
transform 1 0 1308 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_14
timestamp 1714281807
transform 1 0 1212 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_15
timestamp 1714281807
transform 1 0 1252 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_16
timestamp 1714281807
transform 1 0 1148 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_17
timestamp 1714281807
transform 1 0 1100 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_18
timestamp 1714281807
transform 1 0 996 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_19
timestamp 1714281807
transform 1 0 468 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_20
timestamp 1714281807
transform 1 0 412 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_21
timestamp 1714281807
transform 1 0 332 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_22
timestamp 1714281807
transform 1 0 284 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_23
timestamp 1714281807
transform 1 0 2124 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_24
timestamp 1714281807
transform 1 0 2052 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_25
timestamp 1714281807
transform 1 0 1668 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_26
timestamp 1714281807
transform 1 0 2052 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_27
timestamp 1714281807
transform 1 0 1724 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_28
timestamp 1714281807
transform 1 0 1620 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_29
timestamp 1714281807
transform 1 0 1996 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_30
timestamp 1714281807
transform 1 0 1900 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_31
timestamp 1714281807
transform 1 0 1852 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_32
timestamp 1714281807
transform 1 0 1740 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_33
timestamp 1714281807
transform 1 0 1972 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_34
timestamp 1714281807
transform 1 0 1860 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_35
timestamp 1714281807
transform 1 0 1812 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_36
timestamp 1714281807
transform 1 0 2028 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_37
timestamp 1714281807
transform 1 0 1932 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_38
timestamp 1714281807
transform 1 0 1652 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_39
timestamp 1714281807
transform 1 0 2036 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_40
timestamp 1714281807
transform 1 0 1988 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_41
timestamp 1714281807
transform 1 0 1980 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_42
timestamp 1714281807
transform 1 0 1772 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_43
timestamp 1714281807
transform 1 0 1412 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_44
timestamp 1714281807
transform 1 0 1292 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_45
timestamp 1714281807
transform 1 0 1180 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_46
timestamp 1714281807
transform 1 0 1332 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_47
timestamp 1714281807
transform 1 0 1156 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_48
timestamp 1714281807
transform 1 0 1508 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_49
timestamp 1714281807
transform 1 0 1412 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_50
timestamp 1714281807
transform 1 0 1244 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_51
timestamp 1714281807
transform 1 0 1340 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_52
timestamp 1714281807
transform 1 0 1180 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_53
timestamp 1714281807
transform 1 0 1676 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_54
timestamp 1714281807
transform 1 0 1372 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_55
timestamp 1714281807
transform 1 0 1188 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_56
timestamp 1714281807
transform 1 0 1332 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_57
timestamp 1714281807
transform 1 0 1252 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_58
timestamp 1714281807
transform 1 0 1820 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_59
timestamp 1714281807
transform 1 0 1700 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_60
timestamp 1714281807
transform 1 0 1700 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_61
timestamp 1714281807
transform 1 0 1580 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_62
timestamp 1714281807
transform 1 0 1980 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_63
timestamp 1714281807
transform 1 0 1924 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_64
timestamp 1714281807
transform 1 0 1916 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_65
timestamp 1714281807
transform 1 0 1780 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_66
timestamp 1714281807
transform 1 0 1692 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_67
timestamp 1714281807
transform 1 0 1900 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_68
timestamp 1714281807
transform 1 0 1420 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_69
timestamp 1714281807
transform 1 0 2756 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_70
timestamp 1714281807
transform 1 0 2740 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_71
timestamp 1714281807
transform 1 0 2924 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_72
timestamp 1714281807
transform 1 0 2852 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_73
timestamp 1714281807
transform 1 0 2812 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_74
timestamp 1714281807
transform 1 0 2228 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_75
timestamp 1714281807
transform 1 0 2204 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_76
timestamp 1714281807
transform 1 0 2124 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_77
timestamp 1714281807
transform 1 0 2092 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_78
timestamp 1714281807
transform 1 0 1892 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_79
timestamp 1714281807
transform 1 0 1844 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_80
timestamp 1714281807
transform 1 0 1772 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_81
timestamp 1714281807
transform 1 0 2644 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_82
timestamp 1714281807
transform 1 0 2540 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_83
timestamp 1714281807
transform 1 0 2356 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_84
timestamp 1714281807
transform 1 0 2260 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_85
timestamp 1714281807
transform 1 0 2476 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_86
timestamp 1714281807
transform 1 0 2412 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_87
timestamp 1714281807
transform 1 0 2292 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_88
timestamp 1714281807
transform 1 0 2292 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_89
timestamp 1714281807
transform 1 0 2484 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_90
timestamp 1714281807
transform 1 0 2444 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_91
timestamp 1714281807
transform 1 0 2300 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_92
timestamp 1714281807
transform 1 0 2276 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_93
timestamp 1714281807
transform 1 0 2428 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_94
timestamp 1714281807
transform 1 0 2428 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_95
timestamp 1714281807
transform 1 0 2220 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_96
timestamp 1714281807
transform 1 0 2220 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_97
timestamp 1714281807
transform 1 0 2900 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_98
timestamp 1714281807
transform 1 0 2796 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_99
timestamp 1714281807
transform 1 0 2620 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_100
timestamp 1714281807
transform 1 0 2524 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_101
timestamp 1714281807
transform 1 0 2900 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_102
timestamp 1714281807
transform 1 0 2748 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_103
timestamp 1714281807
transform 1 0 2844 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_104
timestamp 1714281807
transform 1 0 2748 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_105
timestamp 1714281807
transform 1 0 2724 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_106
timestamp 1714281807
transform 1 0 2548 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_107
timestamp 1714281807
transform 1 0 1556 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_108
timestamp 1714281807
transform 1 0 1460 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_109
timestamp 1714281807
transform 1 0 1396 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_110
timestamp 1714281807
transform 1 0 1628 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_111
timestamp 1714281807
transform 1 0 1580 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_112
timestamp 1714281807
transform 1 0 1548 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_113
timestamp 1714281807
transform 1 0 1540 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_114
timestamp 1714281807
transform 1 0 1524 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_115
timestamp 1714281807
transform 1 0 1420 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_116
timestamp 1714281807
transform 1 0 1564 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_117
timestamp 1714281807
transform 1 0 1548 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_118
timestamp 1714281807
transform 1 0 1524 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_119
timestamp 1714281807
transform 1 0 1468 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_120
timestamp 1714281807
transform 1 0 1468 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_121
timestamp 1714281807
transform 1 0 2020 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_122
timestamp 1714281807
transform 1 0 1940 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_123
timestamp 1714281807
transform 1 0 1924 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_124
timestamp 1714281807
transform 1 0 1924 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_125
timestamp 1714281807
transform 1 0 1908 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_126
timestamp 1714281807
transform 1 0 1828 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_127
timestamp 1714281807
transform 1 0 1828 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_128
timestamp 1714281807
transform 1 0 1804 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_129
timestamp 1714281807
transform 1 0 1836 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_130
timestamp 1714281807
transform 1 0 1724 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_131
timestamp 1714281807
transform 1 0 2164 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_132
timestamp 1714281807
transform 1 0 2060 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_133
timestamp 1714281807
transform 1 0 2772 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_134
timestamp 1714281807
transform 1 0 2708 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_135
timestamp 1714281807
transform 1 0 2764 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_136
timestamp 1714281807
transform 1 0 2724 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_137
timestamp 1714281807
transform 1 0 2700 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_138
timestamp 1714281807
transform 1 0 2700 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_139
timestamp 1714281807
transform 1 0 2676 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_140
timestamp 1714281807
transform 1 0 2484 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_141
timestamp 1714281807
transform 1 0 2292 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_142
timestamp 1714281807
transform 1 0 2356 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_143
timestamp 1714281807
transform 1 0 2204 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_144
timestamp 1714281807
transform 1 0 2092 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_145
timestamp 1714281807
transform 1 0 2380 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_146
timestamp 1714281807
transform 1 0 2284 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_147
timestamp 1714281807
transform 1 0 516 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_148
timestamp 1714281807
transform 1 0 452 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_149
timestamp 1714281807
transform 1 0 980 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_150
timestamp 1714281807
transform 1 0 892 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_151
timestamp 1714281807
transform 1 0 628 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_152
timestamp 1714281807
transform 1 0 812 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_153
timestamp 1714281807
transform 1 0 732 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_154
timestamp 1714281807
transform 1 0 1604 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_155
timestamp 1714281807
transform 1 0 1548 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_156
timestamp 1714281807
transform 1 0 1892 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_157
timestamp 1714281807
transform 1 0 1788 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_158
timestamp 1714281807
transform 1 0 1932 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_159
timestamp 1714281807
transform 1 0 1820 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_160
timestamp 1714281807
transform 1 0 1956 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_161
timestamp 1714281807
transform 1 0 1812 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_162
timestamp 1714281807
transform 1 0 1676 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_163
timestamp 1714281807
transform 1 0 1332 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_164
timestamp 1714281807
transform 1 0 1212 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_165
timestamp 1714281807
transform 1 0 1612 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_166
timestamp 1714281807
transform 1 0 1516 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_167
timestamp 1714281807
transform 1 0 1476 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_168
timestamp 1714281807
transform 1 0 1372 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_169
timestamp 1714281807
transform 1 0 2212 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_170
timestamp 1714281807
transform 1 0 2092 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_171
timestamp 1714281807
transform 1 0 1924 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_172
timestamp 1714281807
transform 1 0 1812 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_173
timestamp 1714281807
transform 1 0 2524 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_174
timestamp 1714281807
transform 1 0 2404 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_175
timestamp 1714281807
transform 1 0 2356 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_176
timestamp 1714281807
transform 1 0 2236 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_177
timestamp 1714281807
transform 1 0 2988 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_178
timestamp 1714281807
transform 1 0 2876 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_179
timestamp 1714281807
transform 1 0 2996 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_180
timestamp 1714281807
transform 1 0 2876 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_181
timestamp 1714281807
transform 1 0 2804 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_182
timestamp 1714281807
transform 1 0 2692 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_183
timestamp 1714281807
transform 1 0 2348 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_184
timestamp 1714281807
transform 1 0 2324 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_185
timestamp 1714281807
transform 1 0 2980 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_186
timestamp 1714281807
transform 1 0 2924 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_187
timestamp 1714281807
transform 1 0 2996 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_188
timestamp 1714281807
transform 1 0 2876 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_189
timestamp 1714281807
transform 1 0 1372 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_190
timestamp 1714281807
transform 1 0 1348 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_191
timestamp 1714281807
transform 1 0 2972 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_192
timestamp 1714281807
transform 1 0 2860 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_193
timestamp 1714281807
transform 1 0 2844 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_194
timestamp 1714281807
transform 1 0 2724 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_195
timestamp 1714281807
transform 1 0 2468 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_196
timestamp 1714281807
transform 1 0 2364 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_197
timestamp 1714281807
transform 1 0 2340 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_198
timestamp 1714281807
transform 1 0 2236 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_199
timestamp 1714281807
transform 1 0 2212 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_200
timestamp 1714281807
transform 1 0 2108 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_201
timestamp 1714281807
transform 1 0 2956 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_202
timestamp 1714281807
transform 1 0 2828 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_203
timestamp 1714281807
transform 1 0 2996 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_204
timestamp 1714281807
transform 1 0 2876 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_205
timestamp 1714281807
transform 1 0 2860 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_206
timestamp 1714281807
transform 1 0 2732 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_207
timestamp 1714281807
transform 1 0 2428 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_208
timestamp 1714281807
transform 1 0 2308 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_209
timestamp 1714281807
transform 1 0 2500 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_210
timestamp 1714281807
transform 1 0 2444 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_211
timestamp 1714281807
transform 1 0 636 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_212
timestamp 1714281807
transform 1 0 580 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_213
timestamp 1714281807
transform 1 0 508 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_214
timestamp 1714281807
transform 1 0 484 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_215
timestamp 1714281807
transform 1 0 436 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_216
timestamp 1714281807
transform 1 0 436 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_217
timestamp 1714281807
transform 1 0 468 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_218
timestamp 1714281807
transform 1 0 332 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_219
timestamp 1714281807
transform 1 0 380 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_220
timestamp 1714281807
transform 1 0 252 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_221
timestamp 1714281807
transform 1 0 284 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_222
timestamp 1714281807
transform 1 0 236 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_223
timestamp 1714281807
transform 1 0 284 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_224
timestamp 1714281807
transform 1 0 260 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_225
timestamp 1714281807
transform 1 0 588 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_226
timestamp 1714281807
transform 1 0 500 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_227
timestamp 1714281807
transform 1 0 892 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_228
timestamp 1714281807
transform 1 0 812 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_229
timestamp 1714281807
transform 1 0 1380 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_230
timestamp 1714281807
transform 1 0 932 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_231
timestamp 1714281807
transform 1 0 884 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_232
timestamp 1714281807
transform 1 0 780 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_233
timestamp 1714281807
transform 1 0 668 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_234
timestamp 1714281807
transform 1 0 660 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_235
timestamp 1714281807
transform 1 0 916 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_236
timestamp 1714281807
transform 1 0 812 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_237
timestamp 1714281807
transform 1 0 1388 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_238
timestamp 1714281807
transform 1 0 1212 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_239
timestamp 1714281807
transform 1 0 1100 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_240
timestamp 1714281807
transform 1 0 1180 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_241
timestamp 1714281807
transform 1 0 1116 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_242
timestamp 1714281807
transform 1 0 1204 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_243
timestamp 1714281807
transform 1 0 1172 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_244
timestamp 1714281807
transform 1 0 1172 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_245
timestamp 1714281807
transform 1 0 1020 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_246
timestamp 1714281807
transform 1 0 1180 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_247
timestamp 1714281807
transform 1 0 1108 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_248
timestamp 1714281807
transform 1 0 940 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_249
timestamp 1714281807
transform 1 0 876 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_250
timestamp 1714281807
transform 1 0 796 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_251
timestamp 1714281807
transform 1 0 636 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_252
timestamp 1714281807
transform 1 0 388 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_253
timestamp 1714281807
transform 1 0 268 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_254
timestamp 1714281807
transform 1 0 444 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_255
timestamp 1714281807
transform 1 0 276 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_256
timestamp 1714281807
transform 1 0 940 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_257
timestamp 1714281807
transform 1 0 836 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_258
timestamp 1714281807
transform 1 0 740 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_259
timestamp 1714281807
transform 1 0 644 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_260
timestamp 1714281807
transform 1 0 548 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_261
timestamp 1714281807
transform 1 0 452 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_262
timestamp 1714281807
transform 1 0 356 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_263
timestamp 1714281807
transform 1 0 964 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_264
timestamp 1714281807
transform 1 0 844 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_265
timestamp 1714281807
transform 1 0 804 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_266
timestamp 1714281807
transform 1 0 700 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_267
timestamp 1714281807
transform 1 0 268 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_268
timestamp 1714281807
transform 1 0 236 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_269
timestamp 1714281807
transform 1 0 228 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_270
timestamp 1714281807
transform 1 0 204 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_271
timestamp 1714281807
transform 1 0 132 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_272
timestamp 1714281807
transform 1 0 132 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_273
timestamp 1714281807
transform 1 0 100 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_274
timestamp 1714281807
transform 1 0 2492 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_275
timestamp 1714281807
transform 1 0 2116 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_276
timestamp 1714281807
transform 1 0 1468 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_277
timestamp 1714281807
transform 1 0 1396 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_278
timestamp 1714281807
transform 1 0 1396 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_279
timestamp 1714281807
transform 1 0 772 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_280
timestamp 1714281807
transform 1 0 772 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_281
timestamp 1714281807
transform 1 0 716 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_282
timestamp 1714281807
transform 1 0 2788 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_283
timestamp 1714281807
transform 1 0 2684 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_284
timestamp 1714281807
transform 1 0 2580 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_285
timestamp 1714281807
transform 1 0 2580 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_286
timestamp 1714281807
transform 1 0 2476 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_287
timestamp 1714281807
transform 1 0 2460 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_288
timestamp 1714281807
transform 1 0 2308 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_289
timestamp 1714281807
transform 1 0 2228 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_290
timestamp 1714281807
transform 1 0 2140 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_291
timestamp 1714281807
transform 1 0 1988 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_292
timestamp 1714281807
transform 1 0 1892 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_293
timestamp 1714281807
transform 1 0 1676 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_294
timestamp 1714281807
transform 1 0 1660 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_295
timestamp 1714281807
transform 1 0 1612 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_296
timestamp 1714281807
transform 1 0 2916 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_297
timestamp 1714281807
transform 1 0 2828 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_298
timestamp 1714281807
transform 1 0 2764 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_299
timestamp 1714281807
transform 1 0 2732 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_300
timestamp 1714281807
transform 1 0 2628 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_301
timestamp 1714281807
transform 1 0 2628 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_302
timestamp 1714281807
transform 1 0 2628 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_303
timestamp 1714281807
transform 1 0 2596 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_304
timestamp 1714281807
transform 1 0 2500 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_305
timestamp 1714281807
transform 1 0 2484 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_306
timestamp 1714281807
transform 1 0 2484 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_307
timestamp 1714281807
transform 1 0 2412 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_308
timestamp 1714281807
transform 1 0 2404 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_309
timestamp 1714281807
transform 1 0 2308 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_310
timestamp 1714281807
transform 1 0 2132 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_311
timestamp 1714281807
transform 1 0 2108 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_312
timestamp 1714281807
transform 1 0 1900 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_313
timestamp 1714281807
transform 1 0 1748 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_314
timestamp 1714281807
transform 1 0 1740 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_315
timestamp 1714281807
transform 1 0 1636 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_316
timestamp 1714281807
transform 1 0 1636 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_317
timestamp 1714281807
transform 1 0 1588 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_318
timestamp 1714281807
transform 1 0 1428 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_319
timestamp 1714281807
transform 1 0 1252 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_320
timestamp 1714281807
transform 1 0 1076 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_321
timestamp 1714281807
transform 1 0 1052 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_322
timestamp 1714281807
transform 1 0 956 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_323
timestamp 1714281807
transform 1 0 956 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_324
timestamp 1714281807
transform 1 0 2980 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_325
timestamp 1714281807
transform 1 0 2980 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_326
timestamp 1714281807
transform 1 0 2884 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_327
timestamp 1714281807
transform 1 0 2876 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_328
timestamp 1714281807
transform 1 0 2356 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_329
timestamp 1714281807
transform 1 0 2244 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_330
timestamp 1714281807
transform 1 0 2236 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_331
timestamp 1714281807
transform 1 0 2148 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_332
timestamp 1714281807
transform 1 0 2132 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_333
timestamp 1714281807
transform 1 0 2084 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_334
timestamp 1714281807
transform 1 0 1996 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_335
timestamp 1714281807
transform 1 0 1748 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_336
timestamp 1714281807
transform 1 0 1724 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_337
timestamp 1714281807
transform 1 0 1724 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_338
timestamp 1714281807
transform 1 0 1620 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_339
timestamp 1714281807
transform 1 0 1588 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_340
timestamp 1714281807
transform 1 0 2964 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_341
timestamp 1714281807
transform 1 0 2964 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_342
timestamp 1714281807
transform 1 0 2884 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_343
timestamp 1714281807
transform 1 0 2876 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_344
timestamp 1714281807
transform 1 0 2828 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_345
timestamp 1714281807
transform 1 0 2788 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_346
timestamp 1714281807
transform 1 0 2540 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_347
timestamp 1714281807
transform 1 0 2540 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_348
timestamp 1714281807
transform 1 0 2476 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_349
timestamp 1714281807
transform 1 0 2476 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_350
timestamp 1714281807
transform 1 0 2300 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_351
timestamp 1714281807
transform 1 0 2292 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_352
timestamp 1714281807
transform 1 0 2004 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_353
timestamp 1714281807
transform 1 0 2004 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_354
timestamp 1714281807
transform 1 0 1756 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_355
timestamp 1714281807
transform 1 0 1740 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_356
timestamp 1714281807
transform 1 0 1660 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_357
timestamp 1714281807
transform 1 0 2868 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_358
timestamp 1714281807
transform 1 0 2788 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_359
timestamp 1714281807
transform 1 0 2588 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_360
timestamp 1714281807
transform 1 0 2580 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_361
timestamp 1714281807
transform 1 0 2548 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_362
timestamp 1714281807
transform 1 0 2356 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_363
timestamp 1714281807
transform 1 0 2356 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_364
timestamp 1714281807
transform 1 0 2172 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_365
timestamp 1714281807
transform 1 0 2124 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_366
timestamp 1714281807
transform 1 0 2084 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_367
timestamp 1714281807
transform 1 0 1836 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_368
timestamp 1714281807
transform 1 0 1572 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_369
timestamp 1714281807
transform 1 0 2180 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_370
timestamp 1714281807
transform 1 0 2092 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_371
timestamp 1714281807
transform 1 0 2076 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_372
timestamp 1714281807
transform 1 0 2076 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_373
timestamp 1714281807
transform 1 0 2036 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_374
timestamp 1714281807
transform 1 0 2020 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_375
timestamp 1714281807
transform 1 0 2020 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_376
timestamp 1714281807
transform 1 0 1868 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_377
timestamp 1714281807
transform 1 0 1668 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_378
timestamp 1714281807
transform 1 0 1548 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_379
timestamp 1714281807
transform 1 0 1524 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_380
timestamp 1714281807
transform 1 0 1524 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_381
timestamp 1714281807
transform 1 0 1516 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_382
timestamp 1714281807
transform 1 0 1476 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_383
timestamp 1714281807
transform 1 0 1412 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_384
timestamp 1714281807
transform 1 0 1300 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_385
timestamp 1714281807
transform 1 0 1188 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_386
timestamp 1714281807
transform 1 0 1116 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_387
timestamp 1714281807
transform 1 0 1076 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_388
timestamp 1714281807
transform 1 0 972 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_389
timestamp 1714281807
transform 1 0 932 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_390
timestamp 1714281807
transform 1 0 884 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_391
timestamp 1714281807
transform 1 0 836 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_392
timestamp 1714281807
transform 1 0 620 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_393
timestamp 1714281807
transform 1 0 516 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_394
timestamp 1714281807
transform 1 0 1020 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_395
timestamp 1714281807
transform 1 0 948 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_396
timestamp 1714281807
transform 1 0 2156 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_397
timestamp 1714281807
transform 1 0 2100 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_398
timestamp 1714281807
transform 1 0 1524 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_399
timestamp 1714281807
transform 1 0 1396 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_400
timestamp 1714281807
transform 1 0 460 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_401
timestamp 1714281807
transform 1 0 460 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_402
timestamp 1714281807
transform 1 0 428 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_403
timestamp 1714281807
transform 1 0 396 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_404
timestamp 1714281807
transform 1 0 876 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_405
timestamp 1714281807
transform 1 0 740 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_406
timestamp 1714281807
transform 1 0 460 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_407
timestamp 1714281807
transform 1 0 1204 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_408
timestamp 1714281807
transform 1 0 1108 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_409
timestamp 1714281807
transform 1 0 1036 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_410
timestamp 1714281807
transform 1 0 1004 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_411
timestamp 1714281807
transform 1 0 884 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_412
timestamp 1714281807
transform 1 0 820 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_413
timestamp 1714281807
transform 1 0 804 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_414
timestamp 1714281807
transform 1 0 740 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_415
timestamp 1714281807
transform 1 0 740 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_416
timestamp 1714281807
transform 1 0 636 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_417
timestamp 1714281807
transform 1 0 540 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_418
timestamp 1714281807
transform 1 0 540 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_419
timestamp 1714281807
transform 1 0 492 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_420
timestamp 1714281807
transform 1 0 484 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_421
timestamp 1714281807
transform 1 0 484 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_422
timestamp 1714281807
transform 1 0 436 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_423
timestamp 1714281807
transform 1 0 68 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_424
timestamp 1714281807
transform 1 0 44 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_425
timestamp 1714281807
transform 1 0 2452 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_426
timestamp 1714281807
transform 1 0 2372 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_427
timestamp 1714281807
transform 1 0 2332 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_428
timestamp 1714281807
transform 1 0 2268 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_429
timestamp 1714281807
transform 1 0 2268 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_430
timestamp 1714281807
transform 1 0 2164 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_431
timestamp 1714281807
transform 1 0 2164 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_432
timestamp 1714281807
transform 1 0 2068 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_433
timestamp 1714281807
transform 1 0 2036 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_434
timestamp 1714281807
transform 1 0 1964 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_435
timestamp 1714281807
transform 1 0 1844 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_436
timestamp 1714281807
transform 1 0 1772 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_437
timestamp 1714281807
transform 1 0 1764 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_438
timestamp 1714281807
transform 1 0 1988 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_439
timestamp 1714281807
transform 1 0 1972 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_440
timestamp 1714281807
transform 1 0 1684 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_441
timestamp 1714281807
transform 1 0 1604 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_442
timestamp 1714281807
transform 1 0 1604 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_443
timestamp 1714281807
transform 1 0 1540 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_444
timestamp 1714281807
transform 1 0 1516 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_445
timestamp 1714281807
transform 1 0 1508 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_446
timestamp 1714281807
transform 1 0 1420 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_447
timestamp 1714281807
transform 1 0 1412 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_448
timestamp 1714281807
transform 1 0 1412 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_449
timestamp 1714281807
transform 1 0 1388 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_450
timestamp 1714281807
transform 1 0 2668 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_451
timestamp 1714281807
transform 1 0 2652 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_452
timestamp 1714281807
transform 1 0 2564 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_453
timestamp 1714281807
transform 1 0 2548 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_454
timestamp 1714281807
transform 1 0 2500 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_455
timestamp 1714281807
transform 1 0 2476 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_456
timestamp 1714281807
transform 1 0 2132 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_457
timestamp 1714281807
transform 1 0 2132 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_458
timestamp 1714281807
transform 1 0 2108 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_459
timestamp 1714281807
transform 1 0 2092 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_460
timestamp 1714281807
transform 1 0 2076 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_461
timestamp 1714281807
transform 1 0 2076 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_462
timestamp 1714281807
transform 1 0 1988 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_463
timestamp 1714281807
transform 1 0 1956 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_464
timestamp 1714281807
transform 1 0 1884 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_465
timestamp 1714281807
transform 1 0 1788 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_466
timestamp 1714281807
transform 1 0 2756 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_467
timestamp 1714281807
transform 1 0 2716 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_468
timestamp 1714281807
transform 1 0 2516 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_469
timestamp 1714281807
transform 1 0 2516 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_470
timestamp 1714281807
transform 1 0 2356 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_471
timestamp 1714281807
transform 1 0 2332 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_472
timestamp 1714281807
transform 1 0 2292 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_473
timestamp 1714281807
transform 1 0 2196 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_474
timestamp 1714281807
transform 1 0 2196 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_475
timestamp 1714281807
transform 1 0 2188 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_476
timestamp 1714281807
transform 1 0 2140 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_477
timestamp 1714281807
transform 1 0 2140 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_478
timestamp 1714281807
transform 1 0 1036 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_479
timestamp 1714281807
transform 1 0 604 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_480
timestamp 1714281807
transform 1 0 1084 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_481
timestamp 1714281807
transform 1 0 1012 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_482
timestamp 1714281807
transform 1 0 316 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_483
timestamp 1714281807
transform 1 0 252 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_484
timestamp 1714281807
transform 1 0 1228 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_485
timestamp 1714281807
transform 1 0 836 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_486
timestamp 1714281807
transform 1 0 820 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_487
timestamp 1714281807
transform 1 0 700 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_488
timestamp 1714281807
transform 1 0 540 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_489
timestamp 1714281807
transform 1 0 1284 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_490
timestamp 1714281807
transform 1 0 1252 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_491
timestamp 1714281807
transform 1 0 1252 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_492
timestamp 1714281807
transform 1 0 1220 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_493
timestamp 1714281807
transform 1 0 1476 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_494
timestamp 1714281807
transform 1 0 1364 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_495
timestamp 1714281807
transform 1 0 1124 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_496
timestamp 1714281807
transform 1 0 1204 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_497
timestamp 1714281807
transform 1 0 1132 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_498
timestamp 1714281807
transform 1 0 684 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_499
timestamp 1714281807
transform 1 0 2844 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_500
timestamp 1714281807
transform 1 0 2820 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_501
timestamp 1714281807
transform 1 0 2788 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_502
timestamp 1714281807
transform 1 0 2732 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_503
timestamp 1714281807
transform 1 0 2724 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_504
timestamp 1714281807
transform 1 0 2724 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_505
timestamp 1714281807
transform 1 0 2572 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_506
timestamp 1714281807
transform 1 0 2572 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_507
timestamp 1714281807
transform 1 0 2572 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_508
timestamp 1714281807
transform 1 0 2556 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_509
timestamp 1714281807
transform 1 0 2556 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_510
timestamp 1714281807
transform 1 0 2516 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_511
timestamp 1714281807
transform 1 0 2396 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_512
timestamp 1714281807
transform 1 0 2348 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_513
timestamp 1714281807
transform 1 0 2348 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_514
timestamp 1714281807
transform 1 0 2220 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_515
timestamp 1714281807
transform 1 0 2212 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_516
timestamp 1714281807
transform 1 0 2204 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_517
timestamp 1714281807
transform 1 0 2108 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_518
timestamp 1714281807
transform 1 0 2108 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_519
timestamp 1714281807
transform 1 0 2092 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_520
timestamp 1714281807
transform 1 0 2068 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_521
timestamp 1714281807
transform 1 0 2020 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_522
timestamp 1714281807
transform 1 0 1996 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_523
timestamp 1714281807
transform 1 0 1988 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_524
timestamp 1714281807
transform 1 0 1988 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_525
timestamp 1714281807
transform 1 0 1956 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_526
timestamp 1714281807
transform 1 0 1956 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_527
timestamp 1714281807
transform 1 0 1844 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_528
timestamp 1714281807
transform 1 0 1708 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_529
timestamp 1714281807
transform 1 0 1676 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_530
timestamp 1714281807
transform 1 0 1596 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_531
timestamp 1714281807
transform 1 0 1508 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_532
timestamp 1714281807
transform 1 0 1500 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_533
timestamp 1714281807
transform 1 0 1500 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_534
timestamp 1714281807
transform 1 0 1348 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_535
timestamp 1714281807
transform 1 0 1236 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_536
timestamp 1714281807
transform 1 0 1188 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_537
timestamp 1714281807
transform 1 0 2852 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_538
timestamp 1714281807
transform 1 0 2836 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_539
timestamp 1714281807
transform 1 0 2820 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_540
timestamp 1714281807
transform 1 0 2796 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_541
timestamp 1714281807
transform 1 0 2780 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_542
timestamp 1714281807
transform 1 0 2724 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_543
timestamp 1714281807
transform 1 0 2684 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_544
timestamp 1714281807
transform 1 0 2636 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_545
timestamp 1714281807
transform 1 0 2580 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_546
timestamp 1714281807
transform 1 0 2572 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_547
timestamp 1714281807
transform 1 0 2508 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_548
timestamp 1714281807
transform 1 0 2500 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_549
timestamp 1714281807
transform 1 0 2500 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_550
timestamp 1714281807
transform 1 0 2492 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_551
timestamp 1714281807
transform 1 0 2492 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_552
timestamp 1714281807
transform 1 0 2468 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_553
timestamp 1714281807
transform 1 0 2460 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_554
timestamp 1714281807
transform 1 0 2460 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_555
timestamp 1714281807
transform 1 0 2420 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_556
timestamp 1714281807
transform 1 0 2420 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_557
timestamp 1714281807
transform 1 0 2396 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_558
timestamp 1714281807
transform 1 0 2388 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_559
timestamp 1714281807
transform 1 0 2284 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_560
timestamp 1714281807
transform 1 0 2268 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_561
timestamp 1714281807
transform 1 0 2260 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_562
timestamp 1714281807
transform 1 0 2252 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_563
timestamp 1714281807
transform 1 0 2236 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_564
timestamp 1714281807
transform 1 0 2092 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_565
timestamp 1714281807
transform 1 0 2076 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_566
timestamp 1714281807
transform 1 0 2060 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_567
timestamp 1714281807
transform 1 0 2052 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_568
timestamp 1714281807
transform 1 0 2028 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_569
timestamp 1714281807
transform 1 0 1612 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_570
timestamp 1714281807
transform 1 0 1588 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_571
timestamp 1714281807
transform 1 0 1548 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_572
timestamp 1714281807
transform 1 0 1468 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_573
timestamp 1714281807
transform 1 0 1452 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_574
timestamp 1714281807
transform 1 0 1060 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_575
timestamp 1714281807
transform 1 0 2668 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_576
timestamp 1714281807
transform 1 0 2628 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_577
timestamp 1714281807
transform 1 0 2564 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_578
timestamp 1714281807
transform 1 0 2460 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_579
timestamp 1714281807
transform 1 0 2460 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_580
timestamp 1714281807
transform 1 0 2412 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_581
timestamp 1714281807
transform 1 0 2412 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_582
timestamp 1714281807
transform 1 0 2404 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_583
timestamp 1714281807
transform 1 0 2228 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_584
timestamp 1714281807
transform 1 0 2076 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_585
timestamp 1714281807
transform 1 0 1964 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_586
timestamp 1714281807
transform 1 0 1948 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_587
timestamp 1714281807
transform 1 0 1804 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_588
timestamp 1714281807
transform 1 0 1308 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_589
timestamp 1714281807
transform 1 0 1068 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_590
timestamp 1714281807
transform 1 0 1036 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_591
timestamp 1714281807
transform 1 0 996 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_592
timestamp 1714281807
transform 1 0 1372 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_593
timestamp 1714281807
transform 1 0 1268 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_594
timestamp 1714281807
transform 1 0 1292 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_595
timestamp 1714281807
transform 1 0 1228 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_596
timestamp 1714281807
transform 1 0 1188 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_597
timestamp 1714281807
transform 1 0 2668 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_598
timestamp 1714281807
transform 1 0 2596 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_599
timestamp 1714281807
transform 1 0 2540 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_600
timestamp 1714281807
transform 1 0 2532 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_601
timestamp 1714281807
transform 1 0 2316 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_602
timestamp 1714281807
transform 1 0 2252 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_603
timestamp 1714281807
transform 1 0 2244 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_604
timestamp 1714281807
transform 1 0 2244 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_605
timestamp 1714281807
transform 1 0 2228 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_606
timestamp 1714281807
transform 1 0 2220 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_607
timestamp 1714281807
transform 1 0 2212 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_608
timestamp 1714281807
transform 1 0 2172 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_609
timestamp 1714281807
transform 1 0 1924 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_610
timestamp 1714281807
transform 1 0 1748 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_611
timestamp 1714281807
transform 1 0 1676 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_612
timestamp 1714281807
transform 1 0 1676 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_613
timestamp 1714281807
transform 1 0 1636 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_614
timestamp 1714281807
transform 1 0 1444 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_615
timestamp 1714281807
transform 1 0 1356 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_616
timestamp 1714281807
transform 1 0 1332 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_617
timestamp 1714281807
transform 1 0 1252 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_618
timestamp 1714281807
transform 1 0 1236 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_619
timestamp 1714281807
transform 1 0 1212 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_620
timestamp 1714281807
transform 1 0 1212 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_621
timestamp 1714281807
transform 1 0 1204 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_622
timestamp 1714281807
transform 1 0 1204 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_623
timestamp 1714281807
transform 1 0 1188 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_624
timestamp 1714281807
transform 1 0 1132 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_625
timestamp 1714281807
transform 1 0 1132 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_626
timestamp 1714281807
transform 1 0 804 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_627
timestamp 1714281807
transform 1 0 732 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_628
timestamp 1714281807
transform 1 0 732 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_629
timestamp 1714281807
transform 1 0 556 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_630
timestamp 1714281807
transform 1 0 396 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_631
timestamp 1714281807
transform 1 0 372 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_632
timestamp 1714281807
transform 1 0 1380 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_633
timestamp 1714281807
transform 1 0 1380 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_634
timestamp 1714281807
transform 1 0 1300 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_635
timestamp 1714281807
transform 1 0 1300 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_636
timestamp 1714281807
transform 1 0 1300 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_637
timestamp 1714281807
transform 1 0 1172 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_638
timestamp 1714281807
transform 1 0 1124 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_639
timestamp 1714281807
transform 1 0 1084 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_640
timestamp 1714281807
transform 1 0 1076 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_641
timestamp 1714281807
transform 1 0 1036 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_642
timestamp 1714281807
transform 1 0 2820 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_643
timestamp 1714281807
transform 1 0 2820 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_644
timestamp 1714281807
transform 1 0 2780 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_645
timestamp 1714281807
transform 1 0 2772 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_646
timestamp 1714281807
transform 1 0 2772 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_647
timestamp 1714281807
transform 1 0 2492 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_648
timestamp 1714281807
transform 1 0 2492 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_649
timestamp 1714281807
transform 1 0 2404 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_650
timestamp 1714281807
transform 1 0 2348 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_651
timestamp 1714281807
transform 1 0 2324 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_652
timestamp 1714281807
transform 1 0 2324 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_653
timestamp 1714281807
transform 1 0 2308 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_654
timestamp 1714281807
transform 1 0 2284 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_655
timestamp 1714281807
transform 1 0 2276 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_656
timestamp 1714281807
transform 1 0 2244 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_657
timestamp 1714281807
transform 1 0 2244 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_658
timestamp 1714281807
transform 1 0 2236 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_659
timestamp 1714281807
transform 1 0 2228 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_660
timestamp 1714281807
transform 1 0 2028 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_661
timestamp 1714281807
transform 1 0 1948 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_662
timestamp 1714281807
transform 1 0 1868 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_663
timestamp 1714281807
transform 1 0 1860 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_664
timestamp 1714281807
transform 1 0 1684 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_665
timestamp 1714281807
transform 1 0 1564 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_666
timestamp 1714281807
transform 1 0 1412 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_667
timestamp 1714281807
transform 1 0 1204 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_668
timestamp 1714281807
transform 1 0 1204 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_669
timestamp 1714281807
transform 1 0 1196 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_670
timestamp 1714281807
transform 1 0 1084 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_671
timestamp 1714281807
transform 1 0 2756 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_672
timestamp 1714281807
transform 1 0 2756 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_673
timestamp 1714281807
transform 1 0 2660 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_674
timestamp 1714281807
transform 1 0 2628 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_675
timestamp 1714281807
transform 1 0 2580 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_676
timestamp 1714281807
transform 1 0 2540 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_677
timestamp 1714281807
transform 1 0 2540 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_678
timestamp 1714281807
transform 1 0 2356 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_679
timestamp 1714281807
transform 1 0 2356 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_680
timestamp 1714281807
transform 1 0 2300 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_681
timestamp 1714281807
transform 1 0 2236 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_682
timestamp 1714281807
transform 1 0 2228 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_683
timestamp 1714281807
transform 1 0 2132 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_684
timestamp 1714281807
transform 1 0 2132 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_685
timestamp 1714281807
transform 1 0 1908 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_686
timestamp 1714281807
transform 1 0 1852 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_687
timestamp 1714281807
transform 1 0 1852 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_688
timestamp 1714281807
transform 1 0 1804 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_689
timestamp 1714281807
transform 1 0 1772 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_690
timestamp 1714281807
transform 1 0 1748 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_691
timestamp 1714281807
transform 1 0 1748 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_692
timestamp 1714281807
transform 1 0 1508 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_693
timestamp 1714281807
transform 1 0 1444 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_694
timestamp 1714281807
transform 1 0 1332 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_695
timestamp 1714281807
transform 1 0 1268 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_696
timestamp 1714281807
transform 1 0 2996 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_697
timestamp 1714281807
transform 1 0 2996 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_698
timestamp 1714281807
transform 1 0 2836 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_699
timestamp 1714281807
transform 1 0 2780 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_700
timestamp 1714281807
transform 1 0 2780 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_701
timestamp 1714281807
transform 1 0 2772 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_702
timestamp 1714281807
transform 1 0 2740 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_703
timestamp 1714281807
transform 1 0 2732 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_704
timestamp 1714281807
transform 1 0 2588 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_705
timestamp 1714281807
transform 1 0 2588 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_706
timestamp 1714281807
transform 1 0 2356 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_707
timestamp 1714281807
transform 1 0 2356 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_708
timestamp 1714281807
transform 1 0 2316 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_709
timestamp 1714281807
transform 1 0 2316 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_710
timestamp 1714281807
transform 1 0 2300 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_711
timestamp 1714281807
transform 1 0 2276 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_712
timestamp 1714281807
transform 1 0 2116 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_713
timestamp 1714281807
transform 1 0 1964 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_714
timestamp 1714281807
transform 1 0 1964 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_715
timestamp 1714281807
transform 1 0 1828 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_716
timestamp 1714281807
transform 1 0 1740 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_717
timestamp 1714281807
transform 1 0 1740 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_718
timestamp 1714281807
transform 1 0 1740 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_719
timestamp 1714281807
transform 1 0 1716 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_720
timestamp 1714281807
transform 1 0 1716 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_721
timestamp 1714281807
transform 1 0 1452 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_722
timestamp 1714281807
transform 1 0 1268 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_723
timestamp 1714281807
transform 1 0 1196 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_724
timestamp 1714281807
transform 1 0 1180 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_725
timestamp 1714281807
transform 1 0 980 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_726
timestamp 1714281807
transform 1 0 972 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_727
timestamp 1714281807
transform 1 0 948 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_728
timestamp 1714281807
transform 1 0 948 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_729
timestamp 1714281807
transform 1 0 884 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_730
timestamp 1714281807
transform 1 0 876 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_731
timestamp 1714281807
transform 1 0 788 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_732
timestamp 1714281807
transform 1 0 564 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_733
timestamp 1714281807
transform 1 0 508 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_734
timestamp 1714281807
transform 1 0 452 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_735
timestamp 1714281807
transform 1 0 444 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_736
timestamp 1714281807
transform 1 0 404 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_737
timestamp 1714281807
transform 1 0 348 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_738
timestamp 1714281807
transform 1 0 340 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_739
timestamp 1714281807
transform 1 0 316 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_740
timestamp 1714281807
transform 1 0 844 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_741
timestamp 1714281807
transform 1 0 788 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_742
timestamp 1714281807
transform 1 0 684 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_743
timestamp 1714281807
transform 1 0 620 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_744
timestamp 1714281807
transform 1 0 620 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_745
timestamp 1714281807
transform 1 0 468 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_746
timestamp 1714281807
transform 1 0 412 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_747
timestamp 1714281807
transform 1 0 1020 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_748
timestamp 1714281807
transform 1 0 892 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_749
timestamp 1714281807
transform 1 0 1212 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_750
timestamp 1714281807
transform 1 0 964 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_751
timestamp 1714281807
transform 1 0 1132 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_752
timestamp 1714281807
transform 1 0 988 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_753
timestamp 1714281807
transform 1 0 1108 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_754
timestamp 1714281807
transform 1 0 1076 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_755
timestamp 1714281807
transform 1 0 1068 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_756
timestamp 1714281807
transform 1 0 948 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_757
timestamp 1714281807
transform 1 0 828 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_758
timestamp 1714281807
transform 1 0 756 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_759
timestamp 1714281807
transform 1 0 732 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_760
timestamp 1714281807
transform 1 0 548 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_761
timestamp 1714281807
transform 1 0 492 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_762
timestamp 1714281807
transform 1 0 428 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_763
timestamp 1714281807
transform 1 0 260 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_764
timestamp 1714281807
transform 1 0 1044 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_765
timestamp 1714281807
transform 1 0 1012 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_766
timestamp 1714281807
transform 1 0 900 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_767
timestamp 1714281807
transform 1 0 1324 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_768
timestamp 1714281807
transform 1 0 1188 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_769
timestamp 1714281807
transform 1 0 1236 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_770
timestamp 1714281807
transform 1 0 1036 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_771
timestamp 1714281807
transform 1 0 1212 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_772
timestamp 1714281807
transform 1 0 1012 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_773
timestamp 1714281807
transform 1 0 516 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_774
timestamp 1714281807
transform 1 0 396 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_775
timestamp 1714281807
transform 1 0 628 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_776
timestamp 1714281807
transform 1 0 380 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_777
timestamp 1714281807
transform 1 0 644 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_778
timestamp 1714281807
transform 1 0 500 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_779
timestamp 1714281807
transform 1 0 996 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_780
timestamp 1714281807
transform 1 0 916 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_781
timestamp 1714281807
transform 1 0 1100 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_782
timestamp 1714281807
transform 1 0 956 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_783
timestamp 1714281807
transform 1 0 1148 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_784
timestamp 1714281807
transform 1 0 1100 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_785
timestamp 1714281807
transform 1 0 972 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_786
timestamp 1714281807
transform 1 0 924 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_787
timestamp 1714281807
transform 1 0 860 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_788
timestamp 1714281807
transform 1 0 1196 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_789
timestamp 1714281807
transform 1 0 1148 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_790
timestamp 1714281807
transform 1 0 1116 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_791
timestamp 1714281807
transform 1 0 372 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_792
timestamp 1714281807
transform 1 0 316 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_793
timestamp 1714281807
transform 1 0 932 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_794
timestamp 1714281807
transform 1 0 796 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_795
timestamp 1714281807
transform 1 0 796 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_796
timestamp 1714281807
transform 1 0 772 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_797
timestamp 1714281807
transform 1 0 796 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_798
timestamp 1714281807
transform 1 0 676 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_799
timestamp 1714281807
transform 1 0 596 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_800
timestamp 1714281807
transform 1 0 852 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_801
timestamp 1714281807
transform 1 0 700 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_802
timestamp 1714281807
transform 1 0 700 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_803
timestamp 1714281807
transform 1 0 548 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_804
timestamp 1714281807
transform 1 0 1100 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_805
timestamp 1714281807
transform 1 0 892 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_806
timestamp 1714281807
transform 1 0 892 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_807
timestamp 1714281807
transform 1 0 828 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_808
timestamp 1714281807
transform 1 0 780 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_809
timestamp 1714281807
transform 1 0 732 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_810
timestamp 1714281807
transform 1 0 724 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_811
timestamp 1714281807
transform 1 0 668 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_812
timestamp 1714281807
transform 1 0 572 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_813
timestamp 1714281807
transform 1 0 540 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_814
timestamp 1714281807
transform 1 0 556 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_815
timestamp 1714281807
transform 1 0 380 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_816
timestamp 1714281807
transform 1 0 676 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_817
timestamp 1714281807
transform 1 0 516 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_818
timestamp 1714281807
transform 1 0 396 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_819
timestamp 1714281807
transform 1 0 308 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_820
timestamp 1714281807
transform 1 0 212 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_821
timestamp 1714281807
transform 1 0 284 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_822
timestamp 1714281807
transform 1 0 236 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_823
timestamp 1714281807
transform 1 0 876 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_824
timestamp 1714281807
transform 1 0 644 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_825
timestamp 1714281807
transform 1 0 972 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_826
timestamp 1714281807
transform 1 0 820 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_827
timestamp 1714281807
transform 1 0 1164 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_828
timestamp 1714281807
transform 1 0 1124 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_829
timestamp 1714281807
transform 1 0 1084 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_830
timestamp 1714281807
transform 1 0 1076 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_831
timestamp 1714281807
transform 1 0 1172 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_832
timestamp 1714281807
transform 1 0 1092 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_833
timestamp 1714281807
transform 1 0 1020 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_834
timestamp 1714281807
transform 1 0 956 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_835
timestamp 1714281807
transform 1 0 468 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_836
timestamp 1714281807
transform 1 0 380 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_837
timestamp 1714281807
transform 1 0 1132 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_838
timestamp 1714281807
transform 1 0 1100 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_839
timestamp 1714281807
transform 1 0 628 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_840
timestamp 1714281807
transform 1 0 580 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_841
timestamp 1714281807
transform 1 0 580 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_842
timestamp 1714281807
transform 1 0 540 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_843
timestamp 1714281807
transform 1 0 540 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_844
timestamp 1714281807
transform 1 0 412 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_845
timestamp 1714281807
transform 1 0 308 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_846
timestamp 1714281807
transform 1 0 308 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_847
timestamp 1714281807
transform 1 0 244 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_848
timestamp 1714281807
transform 1 0 1036 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_849
timestamp 1714281807
transform 1 0 932 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_850
timestamp 1714281807
transform 1 0 812 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_851
timestamp 1714281807
transform 1 0 684 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_852
timestamp 1714281807
transform 1 0 652 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_853
timestamp 1714281807
transform 1 0 532 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_854
timestamp 1714281807
transform 1 0 444 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_855
timestamp 1714281807
transform 1 0 420 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_856
timestamp 1714281807
transform 1 0 420 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_857
timestamp 1714281807
transform 1 0 372 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_858
timestamp 1714281807
transform 1 0 260 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_859
timestamp 1714281807
transform 1 0 204 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_860
timestamp 1714281807
transform 1 0 436 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_861
timestamp 1714281807
transform 1 0 316 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_862
timestamp 1714281807
transform 1 0 932 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_863
timestamp 1714281807
transform 1 0 868 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_864
timestamp 1714281807
transform 1 0 916 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_865
timestamp 1714281807
transform 1 0 764 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_866
timestamp 1714281807
transform 1 0 1044 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_867
timestamp 1714281807
transform 1 0 964 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_868
timestamp 1714281807
transform 1 0 1196 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_869
timestamp 1714281807
transform 1 0 1132 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_870
timestamp 1714281807
transform 1 0 1252 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_871
timestamp 1714281807
transform 1 0 1164 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_872
timestamp 1714281807
transform 1 0 1092 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_873
timestamp 1714281807
transform 1 0 996 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_874
timestamp 1714281807
transform 1 0 628 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_875
timestamp 1714281807
transform 1 0 556 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_876
timestamp 1714281807
transform 1 0 548 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_877
timestamp 1714281807
transform 1 0 492 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_878
timestamp 1714281807
transform 1 0 388 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_879
timestamp 1714281807
transform 1 0 284 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_880
timestamp 1714281807
transform 1 0 524 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_881
timestamp 1714281807
transform 1 0 396 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_882
timestamp 1714281807
transform 1 0 284 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_883
timestamp 1714281807
transform 1 0 212 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_884
timestamp 1714281807
transform 1 0 444 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_885
timestamp 1714281807
transform 1 0 380 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_886
timestamp 1714281807
transform 1 0 268 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_887
timestamp 1714281807
transform 1 0 156 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_888
timestamp 1714281807
transform 1 0 292 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_889
timestamp 1714281807
transform 1 0 180 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_890
timestamp 1714281807
transform 1 0 468 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_891
timestamp 1714281807
transform 1 0 380 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_892
timestamp 1714281807
transform 1 0 676 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_893
timestamp 1714281807
transform 1 0 604 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_894
timestamp 1714281807
transform 1 0 1404 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_895
timestamp 1714281807
transform 1 0 1276 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_896
timestamp 1714281807
transform 1 0 2068 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_897
timestamp 1714281807
transform 1 0 2020 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_898
timestamp 1714281807
transform 1 0 1556 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_899
timestamp 1714281807
transform 1 0 1516 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_900
timestamp 1714281807
transform 1 0 1548 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_901
timestamp 1714281807
transform 1 0 1508 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_902
timestamp 1714281807
transform 1 0 1660 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_903
timestamp 1714281807
transform 1 0 1612 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_904
timestamp 1714281807
transform 1 0 2228 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_905
timestamp 1714281807
transform 1 0 2156 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_906
timestamp 1714281807
transform 1 0 2380 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_907
timestamp 1714281807
transform 1 0 2332 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_908
timestamp 1714281807
transform 1 0 2228 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_909
timestamp 1714281807
transform 1 0 2172 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_910
timestamp 1714281807
transform 1 0 2812 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_911
timestamp 1714281807
transform 1 0 2780 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_912
timestamp 1714281807
transform 1 0 1644 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_913
timestamp 1714281807
transform 1 0 1604 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_914
timestamp 1714281807
transform 1 0 1684 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_915
timestamp 1714281807
transform 1 0 1636 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_916
timestamp 1714281807
transform 1 0 2852 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_917
timestamp 1714281807
transform 1 0 2796 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_918
timestamp 1714281807
transform 1 0 2028 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_919
timestamp 1714281807
transform 1 0 1988 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_920
timestamp 1714281807
transform 1 0 1788 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_921
timestamp 1714281807
transform 1 0 1772 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_922
timestamp 1714281807
transform 1 0 2900 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_923
timestamp 1714281807
transform 1 0 2860 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_924
timestamp 1714281807
transform 1 0 2900 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_925
timestamp 1714281807
transform 1 0 2860 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_926
timestamp 1714281807
transform 1 0 2244 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_927
timestamp 1714281807
transform 1 0 2204 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_928
timestamp 1714281807
transform 1 0 2164 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_929
timestamp 1714281807
transform 1 0 2116 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_930
timestamp 1714281807
transform 1 0 1612 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_931
timestamp 1714281807
transform 1 0 1564 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_932
timestamp 1714281807
transform 1 0 1012 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_933
timestamp 1714281807
transform 1 0 972 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_934
timestamp 1714281807
transform 1 0 1060 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_935
timestamp 1714281807
transform 1 0 964 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_936
timestamp 1714281807
transform 1 0 1012 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_937
timestamp 1714281807
transform 1 0 972 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_938
timestamp 1714281807
transform 1 0 1156 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_939
timestamp 1714281807
transform 1 0 1108 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_940
timestamp 1714281807
transform 1 0 1668 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_941
timestamp 1714281807
transform 1 0 1636 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_942
timestamp 1714281807
transform 1 0 1844 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_943
timestamp 1714281807
transform 1 0 1796 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_944
timestamp 1714281807
transform 1 0 2940 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_945
timestamp 1714281807
transform 1 0 2900 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_946
timestamp 1714281807
transform 1 0 2940 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_947
timestamp 1714281807
transform 1 0 2900 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_948
timestamp 1714281807
transform 1 0 1684 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_949
timestamp 1714281807
transform 1 0 1644 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_950
timestamp 1714281807
transform 1 0 2052 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_951
timestamp 1714281807
transform 1 0 2020 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_952
timestamp 1714281807
transform 1 0 1772 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_953
timestamp 1714281807
transform 1 0 1724 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_954
timestamp 1714281807
transform 1 0 2500 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_955
timestamp 1714281807
transform 1 0 2444 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_956
timestamp 1714281807
transform 1 0 2172 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_957
timestamp 1714281807
transform 1 0 2124 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_958
timestamp 1714281807
transform 1 0 2532 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_959
timestamp 1714281807
transform 1 0 2492 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_960
timestamp 1714281807
transform 1 0 2516 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_961
timestamp 1714281807
transform 1 0 2428 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_962
timestamp 1714281807
transform 1 0 2724 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_963
timestamp 1714281807
transform 1 0 2708 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_964
timestamp 1714281807
transform 1 0 2764 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_965
timestamp 1714281807
transform 1 0 2732 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_966
timestamp 1714281807
transform 1 0 1420 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_967
timestamp 1714281807
transform 1 0 1372 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_968
timestamp 1714281807
transform 1 0 836 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_969
timestamp 1714281807
transform 1 0 796 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_970
timestamp 1714281807
transform 1 0 804 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_971
timestamp 1714281807
transform 1 0 764 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_972
timestamp 1714281807
transform 1 0 348 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_973
timestamp 1714281807
transform 1 0 268 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_974
timestamp 1714281807
transform 1 0 2220 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_975
timestamp 1714281807
transform 1 0 2116 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_976
timestamp 1714281807
transform 1 0 2124 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_977
timestamp 1714281807
transform 1 0 2100 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_978
timestamp 1714281807
transform 1 0 2836 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_979
timestamp 1714281807
transform 1 0 2748 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_980
timestamp 1714281807
transform 1 0 2284 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_981
timestamp 1714281807
transform 1 0 2204 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_982
timestamp 1714281807
transform 1 0 2412 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_983
timestamp 1714281807
transform 1 0 2332 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_984
timestamp 1714281807
transform 1 0 2860 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_985
timestamp 1714281807
transform 1 0 2780 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_986
timestamp 1714281807
transform 1 0 2660 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_987
timestamp 1714281807
transform 1 0 2596 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_988
timestamp 1714281807
transform 1 0 2380 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_989
timestamp 1714281807
transform 1 0 2228 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_990
timestamp 1714281807
transform 1 0 2140 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_991
timestamp 1714281807
transform 1 0 2436 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_992
timestamp 1714281807
transform 1 0 2332 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_993
timestamp 1714281807
transform 1 0 2524 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_994
timestamp 1714281807
transform 1 0 2364 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_995
timestamp 1714281807
transform 1 0 1484 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_996
timestamp 1714281807
transform 1 0 1444 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_997
timestamp 1714281807
transform 1 0 1628 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_998
timestamp 1714281807
transform 1 0 1572 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_999
timestamp 1714281807
transform 1 0 1372 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1000
timestamp 1714281807
transform 1 0 1300 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1001
timestamp 1714281807
transform 1 0 1580 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_1002
timestamp 1714281807
transform 1 0 1508 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_1003
timestamp 1714281807
transform 1 0 1356 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_1004
timestamp 1714281807
transform 1 0 1972 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1005
timestamp 1714281807
transform 1 0 1876 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_1006
timestamp 1714281807
transform 1 0 2036 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1007
timestamp 1714281807
transform 1 0 1972 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1008
timestamp 1714281807
transform 1 0 1956 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1009
timestamp 1714281807
transform 1 0 2692 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1010
timestamp 1714281807
transform 1 0 2636 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1011
timestamp 1714281807
transform 1 0 1804 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1012
timestamp 1714281807
transform 1 0 1764 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1013
timestamp 1714281807
transform 1 0 1916 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_1014
timestamp 1714281807
transform 1 0 1860 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_1015
timestamp 1714281807
transform 1 0 2076 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_1016
timestamp 1714281807
transform 1 0 2028 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_1017
timestamp 1714281807
transform 1 0 1948 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_1018
timestamp 1714281807
transform 1 0 2100 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1019
timestamp 1714281807
transform 1 0 2060 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1020
timestamp 1714281807
transform 1 0 2284 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1021
timestamp 1714281807
transform 1 0 2220 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1022
timestamp 1714281807
transform 1 0 2428 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1023
timestamp 1714281807
transform 1 0 2404 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1024
timestamp 1714281807
transform 1 0 2348 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1025
timestamp 1714281807
transform 1 0 2804 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1026
timestamp 1714281807
transform 1 0 2628 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1027
timestamp 1714281807
transform 1 0 2788 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1028
timestamp 1714281807
transform 1 0 2652 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1029
timestamp 1714281807
transform 1 0 2780 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1030
timestamp 1714281807
transform 1 0 2644 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1031
timestamp 1714281807
transform 1 0 2540 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_1032
timestamp 1714281807
transform 1 0 2476 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_1033
timestamp 1714281807
transform 1 0 2780 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1034
timestamp 1714281807
transform 1 0 2612 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1035
timestamp 1714281807
transform 1 0 2828 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_1036
timestamp 1714281807
transform 1 0 2804 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_1037
timestamp 1714281807
transform 1 0 2692 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_1038
timestamp 1714281807
transform 1 0 2436 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1039
timestamp 1714281807
transform 1 0 2332 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1040
timestamp 1714281807
transform 1 0 2588 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1041
timestamp 1714281807
transform 1 0 2548 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1042
timestamp 1714281807
transform 1 0 2372 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1043
timestamp 1714281807
transform 1 0 2308 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1044
timestamp 1714281807
transform 1 0 2476 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1045
timestamp 1714281807
transform 1 0 2348 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1046
timestamp 1714281807
transform 1 0 2124 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1047
timestamp 1714281807
transform 1 0 2020 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1048
timestamp 1714281807
transform 1 0 2052 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1049
timestamp 1714281807
transform 1 0 1964 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_1050
timestamp 1714281807
transform 1 0 1564 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1051
timestamp 1714281807
transform 1 0 1532 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1052
timestamp 1714281807
transform 1 0 1444 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1053
timestamp 1714281807
transform 1 0 1452 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1054
timestamp 1714281807
transform 1 0 1380 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1055
timestamp 1714281807
transform 1 0 1524 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_1056
timestamp 1714281807
transform 1 0 1500 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_1057
timestamp 1714281807
transform 1 0 1580 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_1058
timestamp 1714281807
transform 1 0 1492 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_1059
timestamp 1714281807
transform 1 0 1428 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_1060
timestamp 1714281807
transform 1 0 1484 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1061
timestamp 1714281807
transform 1 0 1396 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1062
timestamp 1714281807
transform 1 0 1492 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_1063
timestamp 1714281807
transform 1 0 1396 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_1064
timestamp 1714281807
transform 1 0 2052 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1065
timestamp 1714281807
transform 1 0 1964 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1066
timestamp 1714281807
transform 1 0 1860 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1067
timestamp 1714281807
transform 1 0 1780 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1068
timestamp 1714281807
transform 1 0 2220 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1069
timestamp 1714281807
transform 1 0 2172 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1070
timestamp 1714281807
transform 1 0 2092 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1071
timestamp 1714281807
transform 1 0 2124 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1072
timestamp 1714281807
transform 1 0 2020 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1073
timestamp 1714281807
transform 1 0 2540 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1074
timestamp 1714281807
transform 1 0 2476 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1075
timestamp 1714281807
transform 1 0 2572 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1076
timestamp 1714281807
transform 1 0 2508 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1077
timestamp 1714281807
transform 1 0 2404 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1078
timestamp 1714281807
transform 1 0 700 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1079
timestamp 1714281807
transform 1 0 532 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1080
timestamp 1714281807
transform 1 0 612 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_1081
timestamp 1714281807
transform 1 0 516 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_1082
timestamp 1714281807
transform 1 0 908 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1083
timestamp 1714281807
transform 1 0 764 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1084
timestamp 1714281807
transform 1 0 732 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1085
timestamp 1714281807
transform 1 0 676 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1086
timestamp 1714281807
transform 1 0 1004 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1087
timestamp 1714281807
transform 1 0 948 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1088
timestamp 1714281807
transform 1 0 948 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1089
timestamp 1714281807
transform 1 0 932 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1090
timestamp 1714281807
transform 1 0 604 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1091
timestamp 1714281807
transform 1 0 1276 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1092
timestamp 1714281807
transform 1 0 1156 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1093
timestamp 1714281807
transform 1 0 1068 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1094
timestamp 1714281807
transform 1 0 1068 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1095
timestamp 1714281807
transform 1 0 1028 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1096
timestamp 1714281807
transform 1 0 948 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1097
timestamp 1714281807
transform 1 0 1284 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_1098
timestamp 1714281807
transform 1 0 1076 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1099
timestamp 1714281807
transform 1 0 1020 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_1100
timestamp 1714281807
transform 1 0 1004 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1101
timestamp 1714281807
transform 1 0 1284 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1102
timestamp 1714281807
transform 1 0 1220 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1103
timestamp 1714281807
transform 1 0 1164 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1104
timestamp 1714281807
transform 1 0 1156 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1105
timestamp 1714281807
transform 1 0 1316 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1106
timestamp 1714281807
transform 1 0 1100 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1107
timestamp 1714281807
transform 1 0 468 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1108
timestamp 1714281807
transform 1 0 420 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1109
timestamp 1714281807
transform 1 0 1676 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1110
timestamp 1714281807
transform 1 0 1564 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1111
timestamp 1714281807
transform 1 0 1636 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1112
timestamp 1714281807
transform 1 0 1612 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1113
timestamp 1714281807
transform 1 0 1596 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1114
timestamp 1714281807
transform 1 0 1548 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1115
timestamp 1714281807
transform 1 0 1548 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1116
timestamp 1714281807
transform 1 0 1700 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_1117
timestamp 1714281807
transform 1 0 1612 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_1118
timestamp 1714281807
transform 1 0 1372 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_1119
timestamp 1714281807
transform 1 0 1156 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_1120
timestamp 1714281807
transform 1 0 1212 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1121
timestamp 1714281807
transform 1 0 1084 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1122
timestamp 1714281807
transform 1 0 1316 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_1123
timestamp 1714281807
transform 1 0 1180 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_1124
timestamp 1714281807
transform 1 0 1076 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1125
timestamp 1714281807
transform 1 0 1044 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1126
timestamp 1714281807
transform 1 0 1044 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_1127
timestamp 1714281807
transform 1 0 1100 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1128
timestamp 1714281807
transform 1 0 1052 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1129
timestamp 1714281807
transform 1 0 1732 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1130
timestamp 1714281807
transform 1 0 1676 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1131
timestamp 1714281807
transform 1 0 1548 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_1132
timestamp 1714281807
transform 1 0 1540 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1133
timestamp 1714281807
transform 1 0 1500 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1134
timestamp 1714281807
transform 1 0 1500 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_1135
timestamp 1714281807
transform 1 0 1860 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_1136
timestamp 1714281807
transform 1 0 1788 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_1137
timestamp 1714281807
transform 1 0 2132 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1138
timestamp 1714281807
transform 1 0 2084 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1139
timestamp 1714281807
transform 1 0 2036 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1140
timestamp 1714281807
transform 1 0 2084 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1141
timestamp 1714281807
transform 1 0 1972 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1142
timestamp 1714281807
transform 1 0 2276 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1143
timestamp 1714281807
transform 1 0 2276 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_1144
timestamp 1714281807
transform 1 0 2228 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_1145
timestamp 1714281807
transform 1 0 2220 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1146
timestamp 1714281807
transform 1 0 2724 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1147
timestamp 1714281807
transform 1 0 2700 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_1148
timestamp 1714281807
transform 1 0 2332 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_1149
timestamp 1714281807
transform 1 0 2060 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_1150
timestamp 1714281807
transform 1 0 2044 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_1151
timestamp 1714281807
transform 1 0 1956 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1152
timestamp 1714281807
transform 1 0 1956 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_1153
timestamp 1714281807
transform 1 0 1804 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1154
timestamp 1714281807
transform 1 0 1804 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_1155
timestamp 1714281807
transform 1 0 1708 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1156
timestamp 1714281807
transform 1 0 1564 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1157
timestamp 1714281807
transform 1 0 1436 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_1158
timestamp 1714281807
transform 1 0 252 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1159
timestamp 1714281807
transform 1 0 212 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_1160
timestamp 1714281807
transform 1 0 1500 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1161
timestamp 1714281807
transform 1 0 1436 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1162
timestamp 1714281807
transform 1 0 1252 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1163
timestamp 1714281807
transform 1 0 684 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1164
timestamp 1714281807
transform 1 0 868 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1165
timestamp 1714281807
transform 1 0 780 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1166
timestamp 1714281807
transform 1 0 1844 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1167
timestamp 1714281807
transform 1 0 1812 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1168
timestamp 1714281807
transform 1 0 1668 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1169
timestamp 1714281807
transform 1 0 1964 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1170
timestamp 1714281807
transform 1 0 1908 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1171
timestamp 1714281807
transform 1 0 1852 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1172
timestamp 1714281807
transform 1 0 1724 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1173
timestamp 1714281807
transform 1 0 1940 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1174
timestamp 1714281807
transform 1 0 1820 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1175
timestamp 1714281807
transform 1 0 1820 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1176
timestamp 1714281807
transform 1 0 1716 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1177
timestamp 1714281807
transform 1 0 564 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1178
timestamp 1714281807
transform 1 0 540 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1179
timestamp 1714281807
transform 1 0 428 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1180
timestamp 1714281807
transform 1 0 396 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1181
timestamp 1714281807
transform 1 0 1124 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1182
timestamp 1714281807
transform 1 0 1084 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1183
timestamp 1714281807
transform 1 0 1180 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1184
timestamp 1714281807
transform 1 0 1068 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1185
timestamp 1714281807
transform 1 0 772 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1186
timestamp 1714281807
transform 1 0 668 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1187
timestamp 1714281807
transform 1 0 652 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1188
timestamp 1714281807
transform 1 0 748 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1189
timestamp 1714281807
transform 1 0 740 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1190
timestamp 1714281807
transform 1 0 644 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1191
timestamp 1714281807
transform 1 0 636 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1192
timestamp 1714281807
transform 1 0 1132 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_1193
timestamp 1714281807
transform 1 0 796 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_1194
timestamp 1714281807
transform 1 0 1220 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_1195
timestamp 1714281807
transform 1 0 796 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_1196
timestamp 1714281807
transform 1 0 1028 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1197
timestamp 1714281807
transform 1 0 756 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1198
timestamp 1714281807
transform 1 0 1052 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1199
timestamp 1714281807
transform 1 0 788 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1200
timestamp 1714281807
transform 1 0 1396 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_1201
timestamp 1714281807
transform 1 0 1228 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_1202
timestamp 1714281807
transform 1 0 1308 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1203
timestamp 1714281807
transform 1 0 1260 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1204
timestamp 1714281807
transform 1 0 1300 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1205
timestamp 1714281807
transform 1 0 1260 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1206
timestamp 1714281807
transform 1 0 1388 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1207
timestamp 1714281807
transform 1 0 1348 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1208
timestamp 1714281807
transform 1 0 1308 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1209
timestamp 1714281807
transform 1 0 1268 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1210
timestamp 1714281807
transform 1 0 932 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_1211
timestamp 1714281807
transform 1 0 828 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_1212
timestamp 1714281807
transform 1 0 940 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1213
timestamp 1714281807
transform 1 0 908 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1214
timestamp 1714281807
transform 1 0 1004 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_1215
timestamp 1714281807
transform 1 0 956 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_1216
timestamp 1714281807
transform 1 0 852 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1217
timestamp 1714281807
transform 1 0 748 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1218
timestamp 1714281807
transform 1 0 988 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1219
timestamp 1714281807
transform 1 0 956 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1220
timestamp 1714281807
transform 1 0 796 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_1221
timestamp 1714281807
transform 1 0 660 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_1222
timestamp 1714281807
transform 1 0 820 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_1223
timestamp 1714281807
transform 1 0 756 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_1224
timestamp 1714281807
transform 1 0 564 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_1225
timestamp 1714281807
transform 1 0 788 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1226
timestamp 1714281807
transform 1 0 556 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_1227
timestamp 1714281807
transform 1 0 468 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_1228
timestamp 1714281807
transform 1 0 1444 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1229
timestamp 1714281807
transform 1 0 1260 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1230
timestamp 1714281807
transform 1 0 1004 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_1231
timestamp 1714281807
transform 1 0 2220 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1232
timestamp 1714281807
transform 1 0 1468 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1233
timestamp 1714281807
transform 1 0 2236 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1234
timestamp 1714281807
transform 1 0 2204 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1235
timestamp 1714281807
transform 1 0 2380 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1236
timestamp 1714281807
transform 1 0 2220 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1237
timestamp 1714281807
transform 1 0 2404 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1238
timestamp 1714281807
transform 1 0 2356 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1239
timestamp 1714281807
transform 1 0 2468 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1240
timestamp 1714281807
transform 1 0 2364 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1241
timestamp 1714281807
transform 1 0 2764 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1242
timestamp 1714281807
transform 1 0 2540 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1243
timestamp 1714281807
transform 1 0 2876 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_1244
timestamp 1714281807
transform 1 0 2756 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_1245
timestamp 1714281807
transform 1 0 2820 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1246
timestamp 1714281807
transform 1 0 2764 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1247
timestamp 1714281807
transform 1 0 2548 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1248
timestamp 1714281807
transform 1 0 2548 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_1249
timestamp 1714281807
transform 1 0 2428 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1250
timestamp 1714281807
transform 1 0 2412 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_1251
timestamp 1714281807
transform 1 0 2540 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1252
timestamp 1714281807
transform 1 0 2540 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_1253
timestamp 1714281807
transform 1 0 2468 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_1254
timestamp 1714281807
transform 1 0 2444 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1255
timestamp 1714281807
transform 1 0 2412 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_1256
timestamp 1714281807
transform 1 0 1612 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_1257
timestamp 1714281807
transform 1 0 2644 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_1258
timestamp 1714281807
transform 1 0 2500 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_1259
timestamp 1714281807
transform 1 0 2876 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_1260
timestamp 1714281807
transform 1 0 2628 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1261
timestamp 1714281807
transform 1 0 2372 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1262
timestamp 1714281807
transform 1 0 2180 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_1263
timestamp 1714281807
transform 1 0 2244 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1264
timestamp 1714281807
transform 1 0 2188 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1265
timestamp 1714281807
transform 1 0 2020 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_1266
timestamp 1714281807
transform 1 0 1908 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_1267
timestamp 1714281807
transform 1 0 2044 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1268
timestamp 1714281807
transform 1 0 1876 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1269
timestamp 1714281807
transform 1 0 2628 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_1270
timestamp 1714281807
transform 1 0 2292 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_1271
timestamp 1714281807
transform 1 0 2268 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1272
timestamp 1714281807
transform 1 0 2236 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1273
timestamp 1714281807
transform 1 0 2364 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_1274
timestamp 1714281807
transform 1 0 2292 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_1275
timestamp 1714281807
transform 1 0 2700 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1276
timestamp 1714281807
transform 1 0 2620 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1277
timestamp 1714281807
transform 1 0 1460 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_1278
timestamp 1714281807
transform 1 0 1380 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_1279
timestamp 1714281807
transform 1 0 1612 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_1280
timestamp 1714281807
transform 1 0 1476 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_1281
timestamp 1714281807
transform 1 0 1836 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1282
timestamp 1714281807
transform 1 0 1508 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1283
timestamp 1714281807
transform 1 0 2388 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_1284
timestamp 1714281807
transform 1 0 1796 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_1285
timestamp 1714281807
transform 1 0 1732 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_1286
timestamp 1714281807
transform 1 0 1668 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_1287
timestamp 1714281807
transform 1 0 1948 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1288
timestamp 1714281807
transform 1 0 1780 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1289
timestamp 1714281807
transform 1 0 1996 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1290
timestamp 1714281807
transform 1 0 1924 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1291
timestamp 1714281807
transform 1 0 1932 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1292
timestamp 1714281807
transform 1 0 1788 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1293
timestamp 1714281807
transform 1 0 2268 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_1294
timestamp 1714281807
transform 1 0 1940 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_1295
timestamp 1714281807
transform 1 0 1596 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_1296
timestamp 1714281807
transform 1 0 1412 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_1297
timestamp 1714281807
transform 1 0 1812 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1298
timestamp 1714281807
transform 1 0 1612 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1299
timestamp 1714281807
transform 1 0 2676 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_1300
timestamp 1714281807
transform 1 0 2452 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_1301
timestamp 1714281807
transform 1 0 2932 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_1302
timestamp 1714281807
transform 1 0 2668 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_1303
timestamp 1714281807
transform 1 0 2436 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1304
timestamp 1714281807
transform 1 0 2388 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1305
timestamp 1714281807
transform 1 0 2372 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1306
timestamp 1714281807
transform 1 0 2188 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1307
timestamp 1714281807
transform 1 0 2668 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1308
timestamp 1714281807
transform 1 0 2388 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1309
timestamp 1714281807
transform 1 0 1820 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_1310
timestamp 1714281807
transform 1 0 1700 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_1311
timestamp 1714281807
transform 1 0 1764 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1312
timestamp 1714281807
transform 1 0 1764 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1313
timestamp 1714281807
transform 1 0 1724 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1314
timestamp 1714281807
transform 1 0 1708 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1315
timestamp 1714281807
transform 1 0 1652 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1316
timestamp 1714281807
transform 1 0 1420 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1317
timestamp 1714281807
transform 1 0 1860 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1318
timestamp 1714281807
transform 1 0 1636 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1319
timestamp 1714281807
transform 1 0 1396 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_1320
timestamp 1714281807
transform 1 0 1236 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_1321
timestamp 1714281807
transform 1 0 1356 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_1322
timestamp 1714281807
transform 1 0 1204 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_1323
timestamp 1714281807
transform 1 0 1628 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_1324
timestamp 1714281807
transform 1 0 1324 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_1325
timestamp 1714281807
transform 1 0 1420 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_1326
timestamp 1714281807
transform 1 0 932 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_1327
timestamp 1714281807
transform 1 0 940 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_1328
timestamp 1714281807
transform 1 0 836 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_1329
timestamp 1714281807
transform 1 0 724 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1330
timestamp 1714281807
transform 1 0 644 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1331
timestamp 1714281807
transform 1 0 2484 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1332
timestamp 1714281807
transform 1 0 2356 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1333
timestamp 1714281807
transform 1 0 2300 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_1334
timestamp 1714281807
transform 1 0 2300 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1335
timestamp 1714281807
transform 1 0 1508 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_1336
timestamp 1714281807
transform 1 0 2500 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_1337
timestamp 1714281807
transform 1 0 2404 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_1338
timestamp 1714281807
transform 1 0 2364 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_1339
timestamp 1714281807
transform 1 0 2276 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_1340
timestamp 1714281807
transform 1 0 1428 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1341
timestamp 1714281807
transform 1 0 1140 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1342
timestamp 1714281807
transform 1 0 1212 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_1343
timestamp 1714281807
transform 1 0 1044 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_1344
timestamp 1714281807
transform 1 0 1172 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1345
timestamp 1714281807
transform 1 0 1084 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1346
timestamp 1714281807
transform 1 0 1076 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1347
timestamp 1714281807
transform 1 0 1004 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1348
timestamp 1714281807
transform 1 0 1148 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1349
timestamp 1714281807
transform 1 0 756 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1350
timestamp 1714281807
transform 1 0 748 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1351
timestamp 1714281807
transform 1 0 476 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1352
timestamp 1714281807
transform 1 0 2108 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_1353
timestamp 1714281807
transform 1 0 2044 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_1354
timestamp 1714281807
transform 1 0 1940 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_1355
timestamp 1714281807
transform 1 0 1908 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_1356
timestamp 1714281807
transform 1 0 1908 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1357
timestamp 1714281807
transform 1 0 1884 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1358
timestamp 1714281807
transform 1 0 1868 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1359
timestamp 1714281807
transform 1 0 1140 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1360
timestamp 1714281807
transform 1 0 2124 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1361
timestamp 1714281807
transform 1 0 2028 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1362
timestamp 1714281807
transform 1 0 2044 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_1363
timestamp 1714281807
transform 1 0 1956 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_1364
timestamp 1714281807
transform 1 0 1876 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_1365
timestamp 1714281807
transform 1 0 1036 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1366
timestamp 1714281807
transform 1 0 620 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1367
timestamp 1714281807
transform 1 0 620 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1368
timestamp 1714281807
transform 1 0 324 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1369
timestamp 1714281807
transform 1 0 1716 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_1370
timestamp 1714281807
transform 1 0 1660 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1371
timestamp 1714281807
transform 1 0 1660 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_1372
timestamp 1714281807
transform 1 0 1556 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1373
timestamp 1714281807
transform 1 0 1476 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1374
timestamp 1714281807
transform 1 0 1404 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1375
timestamp 1714281807
transform 1 0 1244 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1376
timestamp 1714281807
transform 1 0 1692 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_1377
timestamp 1714281807
transform 1 0 1492 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_1378
timestamp 1714281807
transform 1 0 1412 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_1379
timestamp 1714281807
transform 1 0 1724 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1380
timestamp 1714281807
transform 1 0 1708 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1381
timestamp 1714281807
transform 1 0 1444 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_1382
timestamp 1714281807
transform 1 0 1428 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_1383
timestamp 1714281807
transform 1 0 996 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_1384
timestamp 1714281807
transform 1 0 708 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1385
timestamp 1714281807
transform 1 0 260 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1386
timestamp 1714281807
transform 1 0 1292 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1387
timestamp 1714281807
transform 1 0 1276 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1388
timestamp 1714281807
transform 1 0 1212 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1389
timestamp 1714281807
transform 1 0 1204 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_1390
timestamp 1714281807
transform 1 0 1148 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_1391
timestamp 1714281807
transform 1 0 1068 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1392
timestamp 1714281807
transform 1 0 1060 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_1393
timestamp 1714281807
transform 1 0 1044 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1394
timestamp 1714281807
transform 1 0 1228 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1395
timestamp 1714281807
transform 1 0 1132 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_1396
timestamp 1714281807
transform 1 0 1148 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1397
timestamp 1714281807
transform 1 0 1100 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1398
timestamp 1714281807
transform 1 0 996 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1399
timestamp 1714281807
transform 1 0 764 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_1400
timestamp 1714281807
transform 1 0 484 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_1401
timestamp 1714281807
transform 1 0 252 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_1402
timestamp 1714281807
transform 1 0 1268 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1403
timestamp 1714281807
transform 1 0 1212 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1404
timestamp 1714281807
transform 1 0 1204 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_1405
timestamp 1714281807
transform 1 0 1116 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1406
timestamp 1714281807
transform 1 0 1100 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_1407
timestamp 1714281807
transform 1 0 1236 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1408
timestamp 1714281807
transform 1 0 1172 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1409
timestamp 1714281807
transform 1 0 1092 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1410
timestamp 1714281807
transform 1 0 1012 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1411
timestamp 1714281807
transform 1 0 724 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_1412
timestamp 1714281807
transform 1 0 564 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1413
timestamp 1714281807
transform 1 0 404 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1414
timestamp 1714281807
transform 1 0 1788 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_1415
timestamp 1714281807
transform 1 0 1756 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_1416
timestamp 1714281807
transform 1 0 1620 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_1417
timestamp 1714281807
transform 1 0 1532 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_1418
timestamp 1714281807
transform 1 0 1772 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1419
timestamp 1714281807
transform 1 0 1692 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1420
timestamp 1714281807
transform 1 0 1860 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1421
timestamp 1714281807
transform 1 0 1780 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1422
timestamp 1714281807
transform 1 0 1388 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1423
timestamp 1714281807
transform 1 0 1116 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1424
timestamp 1714281807
transform 1 0 764 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1425
timestamp 1714281807
transform 1 0 620 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1426
timestamp 1714281807
transform 1 0 452 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1427
timestamp 1714281807
transform 1 0 1756 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1428
timestamp 1714281807
transform 1 0 1684 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1429
timestamp 1714281807
transform 1 0 1676 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1430
timestamp 1714281807
transform 1 0 1572 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1431
timestamp 1714281807
transform 1 0 1508 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1432
timestamp 1714281807
transform 1 0 1700 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1433
timestamp 1714281807
transform 1 0 1700 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1434
timestamp 1714281807
transform 1 0 1652 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1435
timestamp 1714281807
transform 1 0 1652 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1436
timestamp 1714281807
transform 1 0 1460 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1437
timestamp 1714281807
transform 1 0 1204 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1438
timestamp 1714281807
transform 1 0 748 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1439
timestamp 1714281807
transform 1 0 588 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1440
timestamp 1714281807
transform 1 0 2428 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1441
timestamp 1714281807
transform 1 0 2380 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1442
timestamp 1714281807
transform 1 0 2340 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1443
timestamp 1714281807
transform 1 0 2260 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1444
timestamp 1714281807
transform 1 0 2260 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1445
timestamp 1714281807
transform 1 0 2244 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_1446
timestamp 1714281807
transform 1 0 1564 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1447
timestamp 1714281807
transform 1 0 2396 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_1448
timestamp 1714281807
transform 1 0 2252 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_1449
timestamp 1714281807
transform 1 0 2444 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1450
timestamp 1714281807
transform 1 0 2340 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1451
timestamp 1714281807
transform 1 0 2436 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1452
timestamp 1714281807
transform 1 0 2332 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1453
timestamp 1714281807
transform 1 0 1476 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1454
timestamp 1714281807
transform 1 0 1284 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1455
timestamp 1714281807
transform 1 0 1316 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1456
timestamp 1714281807
transform 1 0 1252 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1457
timestamp 1714281807
transform 1 0 1036 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1458
timestamp 1714281807
transform 1 0 1196 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1459
timestamp 1714281807
transform 1 0 1116 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1460
timestamp 1714281807
transform 1 0 2860 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1461
timestamp 1714281807
transform 1 0 2828 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1462
timestamp 1714281807
transform 1 0 2764 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1463
timestamp 1714281807
transform 1 0 2764 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1464
timestamp 1714281807
transform 1 0 2692 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1465
timestamp 1714281807
transform 1 0 1492 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1466
timestamp 1714281807
transform 1 0 2868 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1467
timestamp 1714281807
transform 1 0 2764 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1468
timestamp 1714281807
transform 1 0 2788 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1469
timestamp 1714281807
transform 1 0 2724 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1470
timestamp 1714281807
transform 1 0 2772 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1471
timestamp 1714281807
transform 1 0 2732 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1472
timestamp 1714281807
transform 1 0 2900 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1473
timestamp 1714281807
transform 1 0 2820 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1474
timestamp 1714281807
transform 1 0 1436 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1475
timestamp 1714281807
transform 1 0 1372 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1476
timestamp 1714281807
transform 1 0 1316 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1477
timestamp 1714281807
transform 1 0 1156 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1478
timestamp 1714281807
transform 1 0 2428 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1479
timestamp 1714281807
transform 1 0 2396 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1480
timestamp 1714281807
transform 1 0 2308 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1481
timestamp 1714281807
transform 1 0 2220 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_1482
timestamp 1714281807
transform 1 0 2220 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1483
timestamp 1714281807
transform 1 0 2124 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_1484
timestamp 1714281807
transform 1 0 2060 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_1485
timestamp 1714281807
transform 1 0 2052 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_1486
timestamp 1714281807
transform 1 0 1404 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_1487
timestamp 1714281807
transform 1 0 2324 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_1488
timestamp 1714281807
transform 1 0 2228 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_1489
timestamp 1714281807
transform 1 0 2100 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_1490
timestamp 1714281807
transform 1 0 2444 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_1491
timestamp 1714281807
transform 1 0 2388 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_1492
timestamp 1714281807
transform 1 0 1180 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1493
timestamp 1714281807
transform 1 0 1148 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1494
timestamp 1714281807
transform 1 0 1940 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1495
timestamp 1714281807
transform 1 0 1884 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_1496
timestamp 1714281807
transform 1 0 1820 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1497
timestamp 1714281807
transform 1 0 1820 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1498
timestamp 1714281807
transform 1 0 1756 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_1499
timestamp 1714281807
transform 1 0 1740 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1500
timestamp 1714281807
transform 1 0 1660 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1501
timestamp 1714281807
transform 1 0 1396 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1502
timestamp 1714281807
transform 1 0 1900 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_1503
timestamp 1714281807
transform 1 0 1812 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_1504
timestamp 1714281807
transform 1 0 1916 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_1505
timestamp 1714281807
transform 1 0 1756 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_1506
timestamp 1714281807
transform 1 0 1716 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_1507
timestamp 1714281807
transform 1 0 1788 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_1508
timestamp 1714281807
transform 1 0 1732 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_1509
timestamp 1714281807
transform 1 0 1988 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_1510
timestamp 1714281807
transform 1 0 1940 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_1511
timestamp 1714281807
transform 1 0 1324 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1512
timestamp 1714281807
transform 1 0 1300 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1513
timestamp 1714281807
transform 1 0 988 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1514
timestamp 1714281807
transform 1 0 900 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1515
timestamp 1714281807
transform 1 0 2828 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_1516
timestamp 1714281807
transform 1 0 2772 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_1517
timestamp 1714281807
transform 1 0 2692 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_1518
timestamp 1714281807
transform 1 0 2580 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_1519
timestamp 1714281807
transform 1 0 2532 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_1520
timestamp 1714281807
transform 1 0 2524 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1521
timestamp 1714281807
transform 1 0 2508 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_1522
timestamp 1714281807
transform 1 0 1364 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_1523
timestamp 1714281807
transform 1 0 2756 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_1524
timestamp 1714281807
transform 1 0 2716 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_1525
timestamp 1714281807
transform 1 0 2740 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_1526
timestamp 1714281807
transform 1 0 2668 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_1527
timestamp 1714281807
transform 1 0 2596 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_1528
timestamp 1714281807
transform 1 0 2508 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_1529
timestamp 1714281807
transform 1 0 1356 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1530
timestamp 1714281807
transform 1 0 1276 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1531
timestamp 1714281807
transform 1 0 1028 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1532
timestamp 1714281807
transform 1 0 1284 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1533
timestamp 1714281807
transform 1 0 1012 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1534
timestamp 1714281807
transform 1 0 924 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1535
timestamp 1714281807
transform 1 0 1484 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1536
timestamp 1714281807
transform 1 0 1436 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1537
timestamp 1714281807
transform 1 0 1436 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1538
timestamp 1714281807
transform 1 0 1428 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_1539
timestamp 1714281807
transform 1 0 1372 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_1540
timestamp 1714281807
transform 1 0 1348 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1541
timestamp 1714281807
transform 1 0 1252 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1542
timestamp 1714281807
transform 1 0 1428 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_1543
timestamp 1714281807
transform 1 0 1356 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_1544
timestamp 1714281807
transform 1 0 1428 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1545
timestamp 1714281807
transform 1 0 1380 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1546
timestamp 1714281807
transform 1 0 1292 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1547
timestamp 1714281807
transform 1 0 1260 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1548
timestamp 1714281807
transform 1 0 1300 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1549
timestamp 1714281807
transform 1 0 924 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1550
timestamp 1714281807
transform 1 0 796 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1551
timestamp 1714281807
transform 1 0 1012 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1552
timestamp 1714281807
transform 1 0 956 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1553
timestamp 1714281807
transform 1 0 876 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1554
timestamp 1714281807
transform 1 0 452 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1555
timestamp 1714281807
transform 1 0 452 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1556
timestamp 1714281807
transform 1 0 420 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1557
timestamp 1714281807
transform 1 0 348 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1558
timestamp 1714281807
transform 1 0 2764 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_1559
timestamp 1714281807
transform 1 0 2556 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1560
timestamp 1714281807
transform 1 0 2556 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_1561
timestamp 1714281807
transform 1 0 1372 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1562
timestamp 1714281807
transform 1 0 2852 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_1563
timestamp 1714281807
transform 1 0 2756 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_1564
timestamp 1714281807
transform 1 0 2700 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_1565
timestamp 1714281807
transform 1 0 2572 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_1566
timestamp 1714281807
transform 1 0 2548 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_1567
timestamp 1714281807
transform 1 0 2652 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1568
timestamp 1714281807
transform 1 0 2564 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1569
timestamp 1714281807
transform 1 0 2860 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1570
timestamp 1714281807
transform 1 0 2756 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_1571
timestamp 1714281807
transform 1 0 1244 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1572
timestamp 1714281807
transform 1 0 1084 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1573
timestamp 1714281807
transform 1 0 1124 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1574
timestamp 1714281807
transform 1 0 1076 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1575
timestamp 1714281807
transform 1 0 892 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1576
timestamp 1714281807
transform 1 0 492 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1577
timestamp 1714281807
transform 1 0 492 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_1578
timestamp 1714281807
transform 1 0 404 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_1579
timestamp 1714281807
transform 1 0 292 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_1580
timestamp 1714281807
transform 1 0 2284 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1581
timestamp 1714281807
transform 1 0 2220 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1582
timestamp 1714281807
transform 1 0 2204 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1583
timestamp 1714281807
transform 1 0 2196 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1584
timestamp 1714281807
transform 1 0 2148 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1585
timestamp 1714281807
transform 1 0 1484 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1586
timestamp 1714281807
transform 1 0 2364 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1587
timestamp 1714281807
transform 1 0 2300 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_1588
timestamp 1714281807
transform 1 0 2348 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_1589
timestamp 1714281807
transform 1 0 2300 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_1590
timestamp 1714281807
transform 1 0 1444 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_1591
timestamp 1714281807
transform 1 0 1284 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1592
timestamp 1714281807
transform 1 0 1188 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1593
timestamp 1714281807
transform 1 0 980 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1594
timestamp 1714281807
transform 1 0 868 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1595
timestamp 1714281807
transform 1 0 1140 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1596
timestamp 1714281807
transform 1 0 1060 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1597
timestamp 1714281807
transform 1 0 908 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1598
timestamp 1714281807
transform 1 0 908 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1599
timestamp 1714281807
transform 1 0 548 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1600
timestamp 1714281807
transform 1 0 508 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1601
timestamp 1714281807
transform 1 0 260 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1602
timestamp 1714281807
transform 1 0 2820 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1603
timestamp 1714281807
transform 1 0 2764 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1604
timestamp 1714281807
transform 1 0 2748 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1605
timestamp 1714281807
transform 1 0 2620 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1606
timestamp 1714281807
transform 1 0 1772 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_1607
timestamp 1714281807
transform 1 0 1764 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1608
timestamp 1714281807
transform 1 0 1428 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_1609
timestamp 1714281807
transform 1 0 2764 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_1610
timestamp 1714281807
transform 1 0 2724 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_1611
timestamp 1714281807
transform 1 0 2692 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1612
timestamp 1714281807
transform 1 0 2660 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1613
timestamp 1714281807
transform 1 0 940 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_1614
timestamp 1714281807
transform 1 0 852 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_1615
timestamp 1714281807
transform 1 0 956 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1616
timestamp 1714281807
transform 1 0 948 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1617
timestamp 1714281807
transform 1 0 924 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1618
timestamp 1714281807
transform 1 0 828 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1619
timestamp 1714281807
transform 1 0 828 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1620
timestamp 1714281807
transform 1 0 2860 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_1621
timestamp 1714281807
transform 1 0 2764 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_1622
timestamp 1714281807
transform 1 0 1388 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1623
timestamp 1714281807
transform 1 0 1236 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1624
timestamp 1714281807
transform 1 0 1244 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1625
timestamp 1714281807
transform 1 0 692 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1626
timestamp 1714281807
transform 1 0 676 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1627
timestamp 1714281807
transform 1 0 620 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1628
timestamp 1714281807
transform 1 0 1260 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1629
timestamp 1714281807
transform 1 0 1220 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_1630
timestamp 1714281807
transform 1 0 1188 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_1631
timestamp 1714281807
transform 1 0 860 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1632
timestamp 1714281807
transform 1 0 860 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1633
timestamp 1714281807
transform 1 0 700 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1634
timestamp 1714281807
transform 1 0 300 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1635
timestamp 1714281807
transform 1 0 292 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_1636
timestamp 1714281807
transform 1 0 268 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_1637
timestamp 1714281807
transform 1 0 268 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1638
timestamp 1714281807
transform 1 0 244 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1639
timestamp 1714281807
transform 1 0 892 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1640
timestamp 1714281807
transform 1 0 804 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1641
timestamp 1714281807
transform 1 0 492 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1642
timestamp 1714281807
transform 1 0 484 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1643
timestamp 1714281807
transform 1 0 420 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_1644
timestamp 1714281807
transform 1 0 404 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1645
timestamp 1714281807
transform 1 0 740 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1646
timestamp 1714281807
transform 1 0 436 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1647
timestamp 1714281807
transform 1 0 1036 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1648
timestamp 1714281807
transform 1 0 860 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1649
timestamp 1714281807
transform 1 0 964 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1650
timestamp 1714281807
transform 1 0 868 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1651
timestamp 1714281807
transform 1 0 948 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_1652
timestamp 1714281807
transform 1 0 900 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_1653
timestamp 1714281807
transform 1 0 1108 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1654
timestamp 1714281807
transform 1 0 1036 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1655
timestamp 1714281807
transform 1 0 564 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_1656
timestamp 1714281807
transform 1 0 428 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_1657
timestamp 1714281807
transform 1 0 604 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1658
timestamp 1714281807
transform 1 0 532 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1659
timestamp 1714281807
transform 1 0 548 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_1660
timestamp 1714281807
transform 1 0 484 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_1661
timestamp 1714281807
transform 1 0 444 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_1662
timestamp 1714281807
transform 1 0 708 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1663
timestamp 1714281807
transform 1 0 620 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1664
timestamp 1714281807
transform 1 0 532 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1665
timestamp 1714281807
transform 1 0 468 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1666
timestamp 1714281807
transform 1 0 692 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1667
timestamp 1714281807
transform 1 0 588 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1668
timestamp 1714281807
transform 1 0 564 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1669
timestamp 1714281807
transform 1 0 532 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1670
timestamp 1714281807
transform 1 0 612 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1671
timestamp 1714281807
transform 1 0 548 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1672
timestamp 1714281807
transform 1 0 484 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1673
timestamp 1714281807
transform 1 0 2116 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1674
timestamp 1714281807
transform 1 0 2020 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1675
timestamp 1714281807
transform 1 0 2780 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_1676
timestamp 1714281807
transform 1 0 2732 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_1677
timestamp 1714281807
transform 1 0 2444 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1678
timestamp 1714281807
transform 1 0 2444 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_1679
timestamp 1714281807
transform 1 0 2068 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1680
timestamp 1714281807
transform 1 0 2052 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1681
timestamp 1714281807
transform 1 0 3076 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1682
timestamp 1714281807
transform 1 0 3036 0 1 25
box -3 -3 3 3
use M3_M2  M3_M2_1683
timestamp 1714281807
transform 1 0 2956 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_1684
timestamp 1714281807
transform 1 0 2956 0 1 25
box -3 -3 3 3
use M3_M2  M3_M2_1685
timestamp 1714281807
transform 1 0 2772 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1686
timestamp 1714281807
transform 1 0 2772 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_1687
timestamp 1714281807
transform 1 0 2740 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1688
timestamp 1714281807
transform 1 0 2468 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1689
timestamp 1714281807
transform 1 0 2028 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1690
timestamp 1714281807
transform 1 0 1900 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1691
timestamp 1714281807
transform 1 0 2964 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1692
timestamp 1714281807
transform 1 0 2964 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_1693
timestamp 1714281807
transform 1 0 2660 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_1694
timestamp 1714281807
transform 1 0 2660 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_1695
timestamp 1714281807
transform 1 0 2444 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_1696
timestamp 1714281807
transform 1 0 2372 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_1697
timestamp 1714281807
transform 1 0 2188 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1698
timestamp 1714281807
transform 1 0 2188 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_1699
timestamp 1714281807
transform 1 0 1956 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1700
timestamp 1714281807
transform 1 0 2668 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1701
timestamp 1714281807
transform 1 0 2492 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_1702
timestamp 1714281807
transform 1 0 2252 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1703
timestamp 1714281807
transform 1 0 2252 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1704
timestamp 1714281807
transform 1 0 2244 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_1705
timestamp 1714281807
transform 1 0 2164 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1706
timestamp 1714281807
transform 1 0 2108 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1707
timestamp 1714281807
transform 1 0 2060 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1708
timestamp 1714281807
transform 1 0 2060 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1709
timestamp 1714281807
transform 1 0 2020 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1710
timestamp 1714281807
transform 1 0 2484 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1711
timestamp 1714281807
transform 1 0 2484 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_1712
timestamp 1714281807
transform 1 0 2340 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_1713
timestamp 1714281807
transform 1 0 2164 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_1714
timestamp 1714281807
transform 1 0 2020 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1715
timestamp 1714281807
transform 1 0 2020 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1716
timestamp 1714281807
transform 1 0 1948 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_1717
timestamp 1714281807
transform 1 0 1948 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1718
timestamp 1714281807
transform 1 0 1836 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_1719
timestamp 1714281807
transform 1 0 2044 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_1720
timestamp 1714281807
transform 1 0 1980 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_1721
timestamp 1714281807
transform 1 0 1444 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1722
timestamp 1714281807
transform 1 0 1428 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_1723
timestamp 1714281807
transform 1 0 652 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1724
timestamp 1714281807
transform 1 0 652 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_1725
timestamp 1714281807
transform 1 0 292 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_1726
timestamp 1714281807
transform 1 0 260 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_1727
timestamp 1714281807
transform 1 0 2108 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1728
timestamp 1714281807
transform 1 0 1924 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_1729
timestamp 1714281807
transform 1 0 1900 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_1730
timestamp 1714281807
transform 1 0 1764 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1731
timestamp 1714281807
transform 1 0 1572 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_1732
timestamp 1714281807
transform 1 0 1572 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_1733
timestamp 1714281807
transform 1 0 68 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_1734
timestamp 1714281807
transform 1 0 68 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1735
timestamp 1714281807
transform 1 0 2948 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1736
timestamp 1714281807
transform 1 0 2948 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1737
timestamp 1714281807
transform 1 0 2716 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_1738
timestamp 1714281807
transform 1 0 2364 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_1739
timestamp 1714281807
transform 1 0 2340 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_1740
timestamp 1714281807
transform 1 0 2028 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_1741
timestamp 1714281807
transform 1 0 1788 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_1742
timestamp 1714281807
transform 1 0 1780 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_1743
timestamp 1714281807
transform 1 0 1500 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_1744
timestamp 1714281807
transform 1 0 2988 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_1745
timestamp 1714281807
transform 1 0 2988 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_1746
timestamp 1714281807
transform 1 0 2620 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_1747
timestamp 1714281807
transform 1 0 2260 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_1748
timestamp 1714281807
transform 1 0 2172 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_1749
timestamp 1714281807
transform 1 0 2172 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1750
timestamp 1714281807
transform 1 0 1988 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_1751
timestamp 1714281807
transform 1 0 1700 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1752
timestamp 1714281807
transform 1 0 1420 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_1753
timestamp 1714281807
transform 1 0 2500 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_1754
timestamp 1714281807
transform 1 0 2140 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_1755
timestamp 1714281807
transform 1 0 2140 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1756
timestamp 1714281807
transform 1 0 1892 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1757
timestamp 1714281807
transform 1 0 1868 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1758
timestamp 1714281807
transform 1 0 1868 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1759
timestamp 1714281807
transform 1 0 1564 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1760
timestamp 1714281807
transform 1 0 1556 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_1761
timestamp 1714281807
transform 1 0 2044 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1762
timestamp 1714281807
transform 1 0 2004 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1763
timestamp 1714281807
transform 1 0 1932 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1764
timestamp 1714281807
transform 1 0 1956 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_1765
timestamp 1714281807
transform 1 0 1916 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_1766
timestamp 1714281807
transform 1 0 2036 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_1767
timestamp 1714281807
transform 1 0 1972 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_1768
timestamp 1714281807
transform 1 0 1860 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_1769
timestamp 1714281807
transform 1 0 1828 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_1770
timestamp 1714281807
transform 1 0 1740 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_1771
timestamp 1714281807
transform 1 0 1980 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1772
timestamp 1714281807
transform 1 0 1972 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1773
timestamp 1714281807
transform 1 0 1972 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_1774
timestamp 1714281807
transform 1 0 1940 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1775
timestamp 1714281807
transform 1 0 1924 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1776
timestamp 1714281807
transform 1 0 1884 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1777
timestamp 1714281807
transform 1 0 1820 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1778
timestamp 1714281807
transform 1 0 1804 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1779
timestamp 1714281807
transform 1 0 1644 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1780
timestamp 1714281807
transform 1 0 1580 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1781
timestamp 1714281807
transform 1 0 1516 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1782
timestamp 1714281807
transform 1 0 1316 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_1783
timestamp 1714281807
transform 1 0 1900 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1784
timestamp 1714281807
transform 1 0 1852 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1785
timestamp 1714281807
transform 1 0 1876 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1786
timestamp 1714281807
transform 1 0 1788 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1787
timestamp 1714281807
transform 1 0 1628 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1788
timestamp 1714281807
transform 1 0 1748 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1789
timestamp 1714281807
transform 1 0 1652 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1790
timestamp 1714281807
transform 1 0 1564 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1791
timestamp 1714281807
transform 1 0 1516 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_1792
timestamp 1714281807
transform 1 0 1732 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1793
timestamp 1714281807
transform 1 0 1628 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1794
timestamp 1714281807
transform 1 0 668 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1795
timestamp 1714281807
transform 1 0 324 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1796
timestamp 1714281807
transform 1 0 1204 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_1797
timestamp 1714281807
transform 1 0 1164 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_1798
timestamp 1714281807
transform 1 0 1052 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_1799
timestamp 1714281807
transform 1 0 948 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_1800
timestamp 1714281807
transform 1 0 932 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1801
timestamp 1714281807
transform 1 0 836 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1802
timestamp 1714281807
transform 1 0 700 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1803
timestamp 1714281807
transform 1 0 652 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1804
timestamp 1714281807
transform 1 0 620 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1805
timestamp 1714281807
transform 1 0 604 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_1806
timestamp 1714281807
transform 1 0 516 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_1807
timestamp 1714281807
transform 1 0 476 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_1808
timestamp 1714281807
transform 1 0 396 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_1809
timestamp 1714281807
transform 1 0 420 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_1810
timestamp 1714281807
transform 1 0 316 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_1811
timestamp 1714281807
transform 1 0 228 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1812
timestamp 1714281807
transform 1 0 204 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1813
timestamp 1714281807
transform 1 0 292 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_1814
timestamp 1714281807
transform 1 0 244 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_1815
timestamp 1714281807
transform 1 0 780 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1816
timestamp 1714281807
transform 1 0 740 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1817
timestamp 1714281807
transform 1 0 836 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1818
timestamp 1714281807
transform 1 0 756 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1819
timestamp 1714281807
transform 1 0 420 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1820
timestamp 1714281807
transform 1 0 220 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1821
timestamp 1714281807
transform 1 0 196 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1822
timestamp 1714281807
transform 1 0 492 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1823
timestamp 1714281807
transform 1 0 204 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1824
timestamp 1714281807
transform 1 0 884 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_1825
timestamp 1714281807
transform 1 0 812 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_1826
timestamp 1714281807
transform 1 0 1060 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1827
timestamp 1714281807
transform 1 0 964 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1828
timestamp 1714281807
transform 1 0 1396 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1829
timestamp 1714281807
transform 1 0 1284 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1830
timestamp 1714281807
transform 1 0 740 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1831
timestamp 1714281807
transform 1 0 716 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1832
timestamp 1714281807
transform 1 0 1308 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1833
timestamp 1714281807
transform 1 0 1276 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1834
timestamp 1714281807
transform 1 0 1412 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1835
timestamp 1714281807
transform 1 0 1220 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1836
timestamp 1714281807
transform 1 0 1308 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_1837
timestamp 1714281807
transform 1 0 1260 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_1838
timestamp 1714281807
transform 1 0 1404 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1839
timestamp 1714281807
transform 1 0 1228 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1840
timestamp 1714281807
transform 1 0 1932 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1841
timestamp 1714281807
transform 1 0 1868 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1842
timestamp 1714281807
transform 1 0 1460 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1843
timestamp 1714281807
transform 1 0 1380 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1844
timestamp 1714281807
transform 1 0 1084 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_1845
timestamp 1714281807
transform 1 0 988 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_1846
timestamp 1714281807
transform 1 0 1132 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1847
timestamp 1714281807
transform 1 0 1108 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_1848
timestamp 1714281807
transform 1 0 1124 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1849
timestamp 1714281807
transform 1 0 1028 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1850
timestamp 1714281807
transform 1 0 1108 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_1851
timestamp 1714281807
transform 1 0 1020 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_1852
timestamp 1714281807
transform 1 0 1308 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1853
timestamp 1714281807
transform 1 0 1228 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1854
timestamp 1714281807
transform 1 0 2460 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1855
timestamp 1714281807
transform 1 0 2420 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1856
timestamp 1714281807
transform 1 0 2940 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1857
timestamp 1714281807
transform 1 0 2868 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1858
timestamp 1714281807
transform 1 0 2156 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_1859
timestamp 1714281807
transform 1 0 2092 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_1860
timestamp 1714281807
transform 1 0 1788 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1861
timestamp 1714281807
transform 1 0 1756 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1862
timestamp 1714281807
transform 1 0 2916 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1863
timestamp 1714281807
transform 1 0 2852 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1864
timestamp 1714281807
transform 1 0 1404 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_1865
timestamp 1714281807
transform 1 0 1332 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_1866
timestamp 1714281807
transform 1 0 2940 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_1867
timestamp 1714281807
transform 1 0 2860 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_1868
timestamp 1714281807
transform 1 0 2364 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1869
timestamp 1714281807
transform 1 0 2292 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1870
timestamp 1714281807
transform 1 0 2332 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1871
timestamp 1714281807
transform 1 0 2260 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1872
timestamp 1714281807
transform 1 0 2940 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1873
timestamp 1714281807
transform 1 0 2868 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1874
timestamp 1714281807
transform 1 0 2940 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1875
timestamp 1714281807
transform 1 0 2868 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1876
timestamp 1714281807
transform 1 0 452 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1877
timestamp 1714281807
transform 1 0 372 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1878
timestamp 1714281807
transform 1 0 772 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1879
timestamp 1714281807
transform 1 0 692 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_1880
timestamp 1714281807
transform 1 0 540 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1881
timestamp 1714281807
transform 1 0 396 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1882
timestamp 1714281807
transform 1 0 548 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_1883
timestamp 1714281807
transform 1 0 396 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_1884
timestamp 1714281807
transform 1 0 2468 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1885
timestamp 1714281807
transform 1 0 2364 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1886
timestamp 1714281807
transform 1 0 2380 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1887
timestamp 1714281807
transform 1 0 2308 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1888
timestamp 1714281807
transform 1 0 2044 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1889
timestamp 1714281807
transform 1 0 1980 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_1890
timestamp 1714281807
transform 1 0 1436 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1891
timestamp 1714281807
transform 1 0 1316 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1892
timestamp 1714281807
transform 1 0 1692 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_1893
timestamp 1714281807
transform 1 0 1644 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_1894
timestamp 1714281807
transform 1 0 1444 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1895
timestamp 1714281807
transform 1 0 1308 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_1896
timestamp 1714281807
transform 1 0 1572 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1897
timestamp 1714281807
transform 1 0 1492 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1898
timestamp 1714281807
transform 1 0 1468 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1899
timestamp 1714281807
transform 1 0 1372 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1900
timestamp 1714281807
transform 1 0 1412 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_1901
timestamp 1714281807
transform 1 0 1300 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_1902
timestamp 1714281807
transform 1 0 1556 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1903
timestamp 1714281807
transform 1 0 1476 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_1904
timestamp 1714281807
transform 1 0 2020 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_1905
timestamp 1714281807
transform 1 0 1940 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_1906
timestamp 1714281807
transform 1 0 2020 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1907
timestamp 1714281807
transform 1 0 1948 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1908
timestamp 1714281807
transform 1 0 2156 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1909
timestamp 1714281807
transform 1 0 2076 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1910
timestamp 1714281807
transform 1 0 2108 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1911
timestamp 1714281807
transform 1 0 2020 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1912
timestamp 1714281807
transform 1 0 2004 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1913
timestamp 1714281807
transform 1 0 1964 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1914
timestamp 1714281807
transform 1 0 1988 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_1915
timestamp 1714281807
transform 1 0 1908 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_1916
timestamp 1714281807
transform 1 0 2764 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_1917
timestamp 1714281807
transform 1 0 2700 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_1918
timestamp 1714281807
transform 1 0 2236 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1919
timestamp 1714281807
transform 1 0 2188 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1920
timestamp 1714281807
transform 1 0 468 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1921
timestamp 1714281807
transform 1 0 372 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1922
timestamp 1714281807
transform 1 0 324 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1923
timestamp 1714281807
transform 1 0 284 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1924
timestamp 1714281807
transform 1 0 300 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1925
timestamp 1714281807
transform 1 0 156 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1926
timestamp 1714281807
transform 1 0 340 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1927
timestamp 1714281807
transform 1 0 188 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1928
timestamp 1714281807
transform 1 0 420 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1929
timestamp 1714281807
transform 1 0 324 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1930
timestamp 1714281807
transform 1 0 884 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1931
timestamp 1714281807
transform 1 0 828 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1932
timestamp 1714281807
transform 1 0 1196 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1933
timestamp 1714281807
transform 1 0 1108 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1934
timestamp 1714281807
transform 1 0 1164 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1935
timestamp 1714281807
transform 1 0 1076 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1936
timestamp 1714281807
transform 1 0 2756 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1937
timestamp 1714281807
transform 1 0 2676 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1938
timestamp 1714281807
transform 1 0 2748 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1939
timestamp 1714281807
transform 1 0 2660 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1940
timestamp 1714281807
transform 1 0 2732 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1941
timestamp 1714281807
transform 1 0 2644 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1942
timestamp 1714281807
transform 1 0 604 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1943
timestamp 1714281807
transform 1 0 556 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_1944
timestamp 1714281807
transform 1 0 884 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1945
timestamp 1714281807
transform 1 0 788 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1946
timestamp 1714281807
transform 1 0 764 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1947
timestamp 1714281807
transform 1 0 636 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1948
timestamp 1714281807
transform 1 0 548 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1949
timestamp 1714281807
transform 1 0 780 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1950
timestamp 1714281807
transform 1 0 564 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1951
timestamp 1714281807
transform 1 0 492 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1952
timestamp 1714281807
transform 1 0 676 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_1953
timestamp 1714281807
transform 1 0 572 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_1954
timestamp 1714281807
transform 1 0 548 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1955
timestamp 1714281807
transform 1 0 316 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1956
timestamp 1714281807
transform 1 0 620 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_1957
timestamp 1714281807
transform 1 0 444 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_1958
timestamp 1714281807
transform 1 0 652 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_1959
timestamp 1714281807
transform 1 0 436 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_1960
timestamp 1714281807
transform 1 0 780 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1961
timestamp 1714281807
transform 1 0 692 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1962
timestamp 1714281807
transform 1 0 508 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_1963
timestamp 1714281807
transform 1 0 356 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_1964
timestamp 1714281807
transform 1 0 444 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1965
timestamp 1714281807
transform 1 0 412 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1966
timestamp 1714281807
transform 1 0 788 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_1967
timestamp 1714281807
transform 1 0 508 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_1968
timestamp 1714281807
transform 1 0 516 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1969
timestamp 1714281807
transform 1 0 396 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_1970
timestamp 1714281807
transform 1 0 524 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_1971
timestamp 1714281807
transform 1 0 460 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_1972
timestamp 1714281807
transform 1 0 372 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_1973
timestamp 1714281807
transform 1 0 308 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_1974
timestamp 1714281807
transform 1 0 2052 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1975
timestamp 1714281807
transform 1 0 2004 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1976
timestamp 1714281807
transform 1 0 1996 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_1977
timestamp 1714281807
transform 1 0 1844 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1978
timestamp 1714281807
transform 1 0 1844 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1979
timestamp 1714281807
transform 1 0 1804 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_1980
timestamp 1714281807
transform 1 0 1756 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1981
timestamp 1714281807
transform 1 0 1756 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1982
timestamp 1714281807
transform 1 0 1716 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1983
timestamp 1714281807
transform 1 0 1668 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_1984
timestamp 1714281807
transform 1 0 1668 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1985
timestamp 1714281807
transform 1 0 1668 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_1986
timestamp 1714281807
transform 1 0 1580 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_1987
timestamp 1714281807
transform 1 0 1540 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1988
timestamp 1714281807
transform 1 0 1460 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1989
timestamp 1714281807
transform 1 0 1436 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_1990
timestamp 1714281807
transform 1 0 1436 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1991
timestamp 1714281807
transform 1 0 1076 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1992
timestamp 1714281807
transform 1 0 1044 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1993
timestamp 1714281807
transform 1 0 1036 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1994
timestamp 1714281807
transform 1 0 948 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_1995
timestamp 1714281807
transform 1 0 780 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1996
timestamp 1714281807
transform 1 0 548 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1997
timestamp 1714281807
transform 1 0 828 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_1998
timestamp 1714281807
transform 1 0 740 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_1999
timestamp 1714281807
transform 1 0 892 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_2000
timestamp 1714281807
transform 1 0 668 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_2001
timestamp 1714281807
transform 1 0 892 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2002
timestamp 1714281807
transform 1 0 836 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2003
timestamp 1714281807
transform 1 0 740 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2004
timestamp 1714281807
transform 1 0 508 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2005
timestamp 1714281807
transform 1 0 260 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2006
timestamp 1714281807
transform 1 0 644 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2007
timestamp 1714281807
transform 1 0 516 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2008
timestamp 1714281807
transform 1 0 404 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2009
timestamp 1714281807
transform 1 0 612 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_2010
timestamp 1714281807
transform 1 0 460 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_2011
timestamp 1714281807
transform 1 0 2268 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2012
timestamp 1714281807
transform 1 0 2092 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_2013
timestamp 1714281807
transform 1 0 2204 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_2014
timestamp 1714281807
transform 1 0 2956 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2015
timestamp 1714281807
transform 1 0 2956 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2016
timestamp 1714281807
transform 1 0 3012 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2017
timestamp 1714281807
transform 1 0 2460 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_2018
timestamp 1714281807
transform 1 0 1836 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_2019
timestamp 1714281807
transform 1 0 1836 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_2020
timestamp 1714281807
transform 1 0 1780 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_2021
timestamp 1714281807
transform 1 0 1780 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_2022
timestamp 1714281807
transform 1 0 2956 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_2023
timestamp 1714281807
transform 1 0 2900 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_2024
timestamp 1714281807
transform 1 0 2564 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_2025
timestamp 1714281807
transform 1 0 1740 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2026
timestamp 1714281807
transform 1 0 1740 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_2027
timestamp 1714281807
transform 1 0 1700 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_2028
timestamp 1714281807
transform 1 0 1692 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2029
timestamp 1714281807
transform 1 0 1780 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_2030
timestamp 1714281807
transform 1 0 1772 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_2031
timestamp 1714281807
transform 1 0 1732 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_2032
timestamp 1714281807
transform 1 0 1716 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_2033
timestamp 1714281807
transform 1 0 3012 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_2034
timestamp 1714281807
transform 1 0 2964 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2035
timestamp 1714281807
transform 1 0 2636 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2036
timestamp 1714281807
transform 1 0 2404 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2037
timestamp 1714281807
transform 1 0 2676 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2038
timestamp 1714281807
transform 1 0 2940 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2039
timestamp 1714281807
transform 1 0 2940 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2040
timestamp 1714281807
transform 1 0 2988 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_2041
timestamp 1714281807
transform 1 0 2660 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2042
timestamp 1714281807
transform 1 0 2660 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2043
timestamp 1714281807
transform 1 0 2428 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_2044
timestamp 1714281807
transform 1 0 2308 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2045
timestamp 1714281807
transform 1 0 2252 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2046
timestamp 1714281807
transform 1 0 2340 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2047
timestamp 1714281807
transform 1 0 2340 0 1 75
box -3 -3 3 3
use M3_M2  M3_M2_2048
timestamp 1714281807
transform 1 0 2292 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2049
timestamp 1714281807
transform 1 0 2252 0 1 75
box -3 -3 3 3
use M3_M2  M3_M2_2050
timestamp 1714281807
transform 1 0 2164 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_2051
timestamp 1714281807
transform 1 0 2140 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_2052
timestamp 1714281807
transform 1 0 1748 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2053
timestamp 1714281807
transform 1 0 1748 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2054
timestamp 1714281807
transform 1 0 1684 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2055
timestamp 1714281807
transform 1 0 1684 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2056
timestamp 1714281807
transform 1 0 1612 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2057
timestamp 1714281807
transform 1 0 1604 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_2058
timestamp 1714281807
transform 1 0 1588 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2059
timestamp 1714281807
transform 1 0 1572 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_2060
timestamp 1714281807
transform 1 0 1564 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2061
timestamp 1714281807
transform 1 0 1556 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2062
timestamp 1714281807
transform 1 0 1508 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_2063
timestamp 1714281807
transform 1 0 1508 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2064
timestamp 1714281807
transform 1 0 1716 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_2065
timestamp 1714281807
transform 1 0 1708 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2066
timestamp 1714281807
transform 1 0 1604 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_2067
timestamp 1714281807
transform 1 0 1604 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_2068
timestamp 1714281807
transform 1 0 1500 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2069
timestamp 1714281807
transform 1 0 1468 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_2070
timestamp 1714281807
transform 1 0 2132 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_2071
timestamp 1714281807
transform 1 0 2228 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2072
timestamp 1714281807
transform 1 0 2196 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2073
timestamp 1714281807
transform 1 0 2276 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2074
timestamp 1714281807
transform 1 0 2324 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_2075
timestamp 1714281807
transform 1 0 1956 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2076
timestamp 1714281807
transform 1 0 2596 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_2077
timestamp 1714281807
transform 1 0 2580 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_2078
timestamp 1714281807
transform 1 0 2588 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_2079
timestamp 1714281807
transform 1 0 2644 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_2080
timestamp 1714281807
transform 1 0 2596 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_2081
timestamp 1714281807
transform 1 0 2676 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_2082
timestamp 1714281807
transform 1 0 1684 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_2083
timestamp 1714281807
transform 1 0 1644 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_2084
timestamp 1714281807
transform 1 0 3012 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2085
timestamp 1714281807
transform 1 0 2828 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_2086
timestamp 1714281807
transform 1 0 2676 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2087
timestamp 1714281807
transform 1 0 2580 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2088
timestamp 1714281807
transform 1 0 2572 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2089
timestamp 1714281807
transform 1 0 2740 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2090
timestamp 1714281807
transform 1 0 2988 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2091
timestamp 1714281807
transform 1 0 2988 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2092
timestamp 1714281807
transform 1 0 1020 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2093
timestamp 1714281807
transform 1 0 980 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_2094
timestamp 1714281807
transform 1 0 1156 0 1 55
box -3 -3 3 3
use M3_M2  M3_M2_2095
timestamp 1714281807
transform 1 0 1116 0 1 55
box -3 -3 3 3
use M3_M2  M3_M2_2096
timestamp 1714281807
transform 1 0 2980 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2097
timestamp 1714281807
transform 1 0 2980 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_2098
timestamp 1714281807
transform 1 0 1852 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2099
timestamp 1714281807
transform 1 0 1700 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_2100
timestamp 1714281807
transform 1 0 1676 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_2101
timestamp 1714281807
transform 1 0 1668 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_2102
timestamp 1714281807
transform 1 0 1668 0 1 15
box -3 -3 3 3
use M3_M2  M3_M2_2103
timestamp 1714281807
transform 1 0 140 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_2104
timestamp 1714281807
transform 1 0 140 0 1 15
box -3 -3 3 3
use M3_M2  M3_M2_2105
timestamp 1714281807
transform 1 0 316 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2106
timestamp 1714281807
transform 1 0 348 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_2107
timestamp 1714281807
transform 1 0 292 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_2108
timestamp 1714281807
transform 1 0 236 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_2109
timestamp 1714281807
transform 1 0 324 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2110
timestamp 1714281807
transform 1 0 300 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2111
timestamp 1714281807
transform 1 0 220 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2112
timestamp 1714281807
transform 1 0 172 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_2113
timestamp 1714281807
transform 1 0 796 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2114
timestamp 1714281807
transform 1 0 1524 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_2115
timestamp 1714281807
transform 1 0 1508 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_2116
timestamp 1714281807
transform 1 0 132 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_2117
timestamp 1714281807
transform 1 0 116 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_2118
timestamp 1714281807
transform 1 0 1484 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_2119
timestamp 1714281807
transform 1 0 1452 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2120
timestamp 1714281807
transform 1 0 356 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2121
timestamp 1714281807
transform 1 0 300 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_2122
timestamp 1714281807
transform 1 0 1548 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2123
timestamp 1714281807
transform 1 0 1532 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_2124
timestamp 1714281807
transform 1 0 1500 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2125
timestamp 1714281807
transform 1 0 1500 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_2126
timestamp 1714281807
transform 1 0 1476 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_2127
timestamp 1714281807
transform 1 0 1476 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_2128
timestamp 1714281807
transform 1 0 1452 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_2129
timestamp 1714281807
transform 1 0 1444 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_2130
timestamp 1714281807
transform 1 0 1468 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_2131
timestamp 1714281807
transform 1 0 1468 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_2132
timestamp 1714281807
transform 1 0 1340 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_2133
timestamp 1714281807
transform 1 0 1340 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_2134
timestamp 1714281807
transform 1 0 940 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2135
timestamp 1714281807
transform 1 0 908 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2136
timestamp 1714281807
transform 1 0 916 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2137
timestamp 1714281807
transform 1 0 892 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2138
timestamp 1714281807
transform 1 0 820 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2139
timestamp 1714281807
transform 1 0 732 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2140
timestamp 1714281807
transform 1 0 676 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2141
timestamp 1714281807
transform 1 0 620 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2142
timestamp 1714281807
transform 1 0 532 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2143
timestamp 1714281807
transform 1 0 436 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2144
timestamp 1714281807
transform 1 0 700 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_2145
timestamp 1714281807
transform 1 0 628 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_2146
timestamp 1714281807
transform 1 0 420 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2147
timestamp 1714281807
transform 1 0 1020 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_2148
timestamp 1714281807
transform 1 0 972 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_2149
timestamp 1714281807
transform 1 0 1180 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_2150
timestamp 1714281807
transform 1 0 1164 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_2151
timestamp 1714281807
transform 1 0 1116 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_2152
timestamp 1714281807
transform 1 0 1084 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_2153
timestamp 1714281807
transform 1 0 1060 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_2154
timestamp 1714281807
transform 1 0 1196 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_2155
timestamp 1714281807
transform 1 0 1156 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_2156
timestamp 1714281807
transform 1 0 580 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_2157
timestamp 1714281807
transform 1 0 428 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_2158
timestamp 1714281807
transform 1 0 444 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_2159
timestamp 1714281807
transform 1 0 684 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_2160
timestamp 1714281807
transform 1 0 660 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_2161
timestamp 1714281807
transform 1 0 620 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_2162
timestamp 1714281807
transform 1 0 572 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_2163
timestamp 1714281807
transform 1 0 676 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_2164
timestamp 1714281807
transform 1 0 596 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_2165
timestamp 1714281807
transform 1 0 1556 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2166
timestamp 1714281807
transform 1 0 1556 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_2167
timestamp 1714281807
transform 1 0 1388 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_2168
timestamp 1714281807
transform 1 0 1388 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_2169
timestamp 1714281807
transform 1 0 1732 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_2170
timestamp 1714281807
transform 1 0 1628 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_2171
timestamp 1714281807
transform 1 0 1620 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_2172
timestamp 1714281807
transform 1 0 1620 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_2173
timestamp 1714281807
transform 1 0 1492 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_2174
timestamp 1714281807
transform 1 0 1484 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_2175
timestamp 1714281807
transform 1 0 1428 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_2176
timestamp 1714281807
transform 1 0 1412 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_2177
timestamp 1714281807
transform 1 0 1996 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_2178
timestamp 1714281807
transform 1 0 1932 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_2179
timestamp 1714281807
transform 1 0 1892 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2180
timestamp 1714281807
transform 1 0 1748 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2181
timestamp 1714281807
transform 1 0 1748 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_2182
timestamp 1714281807
transform 1 0 1708 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_2183
timestamp 1714281807
transform 1 0 1708 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2184
timestamp 1714281807
transform 1 0 1636 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_2185
timestamp 1714281807
transform 1 0 1492 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_2186
timestamp 1714281807
transform 1 0 1484 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_2187
timestamp 1714281807
transform 1 0 1316 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_2188
timestamp 1714281807
transform 1 0 1292 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_2189
timestamp 1714281807
transform 1 0 1628 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2190
timestamp 1714281807
transform 1 0 1572 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2191
timestamp 1714281807
transform 1 0 1556 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_2192
timestamp 1714281807
transform 1 0 1508 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_2193
timestamp 1714281807
transform 1 0 1484 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_2194
timestamp 1714281807
transform 1 0 1308 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_2195
timestamp 1714281807
transform 1 0 1276 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_2196
timestamp 1714281807
transform 1 0 892 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_2197
timestamp 1714281807
transform 1 0 860 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2198
timestamp 1714281807
transform 1 0 764 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_2199
timestamp 1714281807
transform 1 0 764 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2200
timestamp 1714281807
transform 1 0 652 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2201
timestamp 1714281807
transform 1 0 628 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2202
timestamp 1714281807
transform 1 0 556 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2203
timestamp 1714281807
transform 1 0 372 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_2204
timestamp 1714281807
transform 1 0 332 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_2205
timestamp 1714281807
transform 1 0 780 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2206
timestamp 1714281807
transform 1 0 628 0 1 85
box -3 -3 3 3
use M3_M2  M3_M2_2207
timestamp 1714281807
transform 1 0 548 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_2208
timestamp 1714281807
transform 1 0 492 0 1 85
box -3 -3 3 3
use M3_M2  M3_M2_2209
timestamp 1714281807
transform 1 0 364 0 1 85
box -3 -3 3 3
use M3_M2  M3_M2_2210
timestamp 1714281807
transform 1 0 348 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2211
timestamp 1714281807
transform 1 0 276 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2212
timestamp 1714281807
transform 1 0 220 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2213
timestamp 1714281807
transform 1 0 588 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_2214
timestamp 1714281807
transform 1 0 476 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_2215
timestamp 1714281807
transform 1 0 324 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_2216
timestamp 1714281807
transform 1 0 772 0 1 75
box -3 -3 3 3
use M3_M2  M3_M2_2217
timestamp 1714281807
transform 1 0 660 0 1 75
box -3 -3 3 3
use M3_M2  M3_M2_2218
timestamp 1714281807
transform 1 0 508 0 1 75
box -3 -3 3 3
use M3_M2  M3_M2_2219
timestamp 1714281807
transform 1 0 380 0 1 75
box -3 -3 3 3
use M3_M2  M3_M2_2220
timestamp 1714281807
transform 1 0 260 0 1 75
box -3 -3 3 3
use M3_M2  M3_M2_2221
timestamp 1714281807
transform 1 0 1012 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2222
timestamp 1714281807
transform 1 0 900 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2223
timestamp 1714281807
transform 1 0 892 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2224
timestamp 1714281807
transform 1 0 844 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2225
timestamp 1714281807
transform 1 0 756 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2226
timestamp 1714281807
transform 1 0 892 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_2227
timestamp 1714281807
transform 1 0 812 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_2228
timestamp 1714281807
transform 1 0 780 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_2229
timestamp 1714281807
transform 1 0 708 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_2230
timestamp 1714281807
transform 1 0 868 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_2231
timestamp 1714281807
transform 1 0 964 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2232
timestamp 1714281807
transform 1 0 948 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_2233
timestamp 1714281807
transform 1 0 716 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_2234
timestamp 1714281807
transform 1 0 508 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_2235
timestamp 1714281807
transform 1 0 452 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_2236
timestamp 1714281807
transform 1 0 172 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_2237
timestamp 1714281807
transform 1 0 172 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2238
timestamp 1714281807
transform 1 0 156 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_2239
timestamp 1714281807
transform 1 0 100 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_2240
timestamp 1714281807
transform 1 0 84 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_2241
timestamp 1714281807
transform 1 0 420 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_2242
timestamp 1714281807
transform 1 0 2036 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_2243
timestamp 1714281807
transform 1 0 1708 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_2244
timestamp 1714281807
transform 1 0 1708 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2245
timestamp 1714281807
transform 1 0 1572 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_2246
timestamp 1714281807
transform 1 0 1476 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2247
timestamp 1714281807
transform 1 0 1404 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2248
timestamp 1714281807
transform 1 0 1404 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_2249
timestamp 1714281807
transform 1 0 1004 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2250
timestamp 1714281807
transform 1 0 2932 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2251
timestamp 1714281807
transform 1 0 2916 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_2252
timestamp 1714281807
transform 1 0 2916 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2253
timestamp 1714281807
transform 1 0 2916 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2254
timestamp 1714281807
transform 1 0 2900 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2255
timestamp 1714281807
transform 1 0 2892 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_2256
timestamp 1714281807
transform 1 0 2868 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_2257
timestamp 1714281807
transform 1 0 2780 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_2258
timestamp 1714281807
transform 1 0 2772 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2259
timestamp 1714281807
transform 1 0 2764 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_2260
timestamp 1714281807
transform 1 0 2764 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_2261
timestamp 1714281807
transform 1 0 2724 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2262
timestamp 1714281807
transform 1 0 2692 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2263
timestamp 1714281807
transform 1 0 2676 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_2264
timestamp 1714281807
transform 1 0 2676 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_2265
timestamp 1714281807
transform 1 0 2676 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2266
timestamp 1714281807
transform 1 0 2676 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2267
timestamp 1714281807
transform 1 0 2668 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2268
timestamp 1714281807
transform 1 0 2652 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2269
timestamp 1714281807
transform 1 0 2628 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_2270
timestamp 1714281807
transform 1 0 2628 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_2271
timestamp 1714281807
transform 1 0 2620 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_2272
timestamp 1714281807
transform 1 0 2612 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2273
timestamp 1714281807
transform 1 0 2612 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2274
timestamp 1714281807
transform 1 0 2612 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_2275
timestamp 1714281807
transform 1 0 2580 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_2276
timestamp 1714281807
transform 1 0 2540 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2277
timestamp 1714281807
transform 1 0 2500 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_2278
timestamp 1714281807
transform 1 0 2492 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_2279
timestamp 1714281807
transform 1 0 2492 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_2280
timestamp 1714281807
transform 1 0 2460 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_2281
timestamp 1714281807
transform 1 0 2444 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_2282
timestamp 1714281807
transform 1 0 2444 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_2283
timestamp 1714281807
transform 1 0 2444 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2284
timestamp 1714281807
transform 1 0 2436 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2285
timestamp 1714281807
transform 1 0 2396 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_2286
timestamp 1714281807
transform 1 0 2388 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_2287
timestamp 1714281807
transform 1 0 2388 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2288
timestamp 1714281807
transform 1 0 2356 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2289
timestamp 1714281807
transform 1 0 2316 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_2290
timestamp 1714281807
transform 1 0 2308 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_2291
timestamp 1714281807
transform 1 0 2308 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2292
timestamp 1714281807
transform 1 0 2276 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2293
timestamp 1714281807
transform 1 0 2268 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2294
timestamp 1714281807
transform 1 0 2260 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_2295
timestamp 1714281807
transform 1 0 2260 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2296
timestamp 1714281807
transform 1 0 2212 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2297
timestamp 1714281807
transform 1 0 2204 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2298
timestamp 1714281807
transform 1 0 2180 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_2299
timestamp 1714281807
transform 1 0 2148 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2300
timestamp 1714281807
transform 1 0 2132 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_2301
timestamp 1714281807
transform 1 0 2132 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2302
timestamp 1714281807
transform 1 0 2124 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2303
timestamp 1714281807
transform 1 0 2124 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2304
timestamp 1714281807
transform 1 0 2124 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2305
timestamp 1714281807
transform 1 0 2116 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2306
timestamp 1714281807
transform 1 0 2084 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_2307
timestamp 1714281807
transform 1 0 2028 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2308
timestamp 1714281807
transform 1 0 2028 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2309
timestamp 1714281807
transform 1 0 1980 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2310
timestamp 1714281807
transform 1 0 1964 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2311
timestamp 1714281807
transform 1 0 1948 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2312
timestamp 1714281807
transform 1 0 1932 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_2313
timestamp 1714281807
transform 1 0 1932 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_2314
timestamp 1714281807
transform 1 0 1916 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2315
timestamp 1714281807
transform 1 0 1900 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2316
timestamp 1714281807
transform 1 0 1900 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_2317
timestamp 1714281807
transform 1 0 1892 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2318
timestamp 1714281807
transform 1 0 1876 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2319
timestamp 1714281807
transform 1 0 1860 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_2320
timestamp 1714281807
transform 1 0 1852 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2321
timestamp 1714281807
transform 1 0 1820 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_2322
timestamp 1714281807
transform 1 0 1820 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2323
timestamp 1714281807
transform 1 0 1812 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2324
timestamp 1714281807
transform 1 0 1812 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2325
timestamp 1714281807
transform 1 0 1804 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2326
timestamp 1714281807
transform 1 0 1756 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_2327
timestamp 1714281807
transform 1 0 1740 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2328
timestamp 1714281807
transform 1 0 1708 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_2329
timestamp 1714281807
transform 1 0 1652 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2330
timestamp 1714281807
transform 1 0 1652 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2331
timestamp 1714281807
transform 1 0 1596 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2332
timestamp 1714281807
transform 1 0 1588 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_2333
timestamp 1714281807
transform 1 0 1588 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2334
timestamp 1714281807
transform 1 0 1532 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2335
timestamp 1714281807
transform 1 0 1524 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_2336
timestamp 1714281807
transform 1 0 1524 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2337
timestamp 1714281807
transform 1 0 1484 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_2338
timestamp 1714281807
transform 1 0 1444 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_2339
timestamp 1714281807
transform 1 0 1428 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2340
timestamp 1714281807
transform 1 0 1404 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_2341
timestamp 1714281807
transform 1 0 1388 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2342
timestamp 1714281807
transform 1 0 1388 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2343
timestamp 1714281807
transform 1 0 1380 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_2344
timestamp 1714281807
transform 1 0 1380 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_2345
timestamp 1714281807
transform 1 0 1332 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2346
timestamp 1714281807
transform 1 0 1308 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_2347
timestamp 1714281807
transform 1 0 1284 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2348
timestamp 1714281807
transform 1 0 1268 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_2349
timestamp 1714281807
transform 1 0 1260 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2350
timestamp 1714281807
transform 1 0 1252 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2351
timestamp 1714281807
transform 1 0 1228 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_2352
timestamp 1714281807
transform 1 0 1172 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_2353
timestamp 1714281807
transform 1 0 1100 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_2354
timestamp 1714281807
transform 1 0 1100 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_2355
timestamp 1714281807
transform 1 0 1068 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2356
timestamp 1714281807
transform 1 0 1068 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2357
timestamp 1714281807
transform 1 0 1060 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_2358
timestamp 1714281807
transform 1 0 1028 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_2359
timestamp 1714281807
transform 1 0 1028 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_2360
timestamp 1714281807
transform 1 0 972 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2361
timestamp 1714281807
transform 1 0 964 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2362
timestamp 1714281807
transform 1 0 948 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_2363
timestamp 1714281807
transform 1 0 948 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_2364
timestamp 1714281807
transform 1 0 852 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_2365
timestamp 1714281807
transform 1 0 836 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2366
timestamp 1714281807
transform 1 0 828 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_2367
timestamp 1714281807
transform 1 0 788 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2368
timestamp 1714281807
transform 1 0 780 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2369
timestamp 1714281807
transform 1 0 772 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2370
timestamp 1714281807
transform 1 0 756 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_2371
timestamp 1714281807
transform 1 0 748 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2372
timestamp 1714281807
transform 1 0 700 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_2373
timestamp 1714281807
transform 1 0 700 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2374
timestamp 1714281807
transform 1 0 604 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_2375
timestamp 1714281807
transform 1 0 572 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2376
timestamp 1714281807
transform 1 0 564 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_2377
timestamp 1714281807
transform 1 0 556 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2378
timestamp 1714281807
transform 1 0 548 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2379
timestamp 1714281807
transform 1 0 508 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2380
timestamp 1714281807
transform 1 0 508 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2381
timestamp 1714281807
transform 1 0 444 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_2382
timestamp 1714281807
transform 1 0 436 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2383
timestamp 1714281807
transform 1 0 436 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2384
timestamp 1714281807
transform 1 0 388 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2385
timestamp 1714281807
transform 1 0 372 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_2386
timestamp 1714281807
transform 1 0 372 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2387
timestamp 1714281807
transform 1 0 364 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2388
timestamp 1714281807
transform 1 0 332 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_2389
timestamp 1714281807
transform 1 0 332 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_2390
timestamp 1714281807
transform 1 0 324 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2391
timestamp 1714281807
transform 1 0 324 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2392
timestamp 1714281807
transform 1 0 308 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2393
timestamp 1714281807
transform 1 0 260 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_2394
timestamp 1714281807
transform 1 0 196 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_2395
timestamp 1714281807
transform 1 0 196 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_2396
timestamp 1714281807
transform 1 0 196 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_2397
timestamp 1714281807
transform 1 0 164 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_2398
timestamp 1714281807
transform 1 0 132 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_2399
timestamp 1714281807
transform 1 0 108 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_2400
timestamp 1714281807
transform 1 0 108 0 1 1185
box -3 -3 3 3
use NAND2X1  NAND2X1_0
timestamp 1714281807
transform 1 0 424 0 1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_1
timestamp 1714281807
transform 1 0 1480 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_2
timestamp 1714281807
transform 1 0 1112 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_3
timestamp 1714281807
transform 1 0 1184 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_4
timestamp 1714281807
transform 1 0 1064 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_5
timestamp 1714281807
transform 1 0 1096 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_6
timestamp 1714281807
transform 1 0 1456 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_7
timestamp 1714281807
transform 1 0 1472 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_8
timestamp 1714281807
transform 1 0 1520 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_9
timestamp 1714281807
transform 1 0 1464 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_10
timestamp 1714281807
transform 1 0 1384 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_11
timestamp 1714281807
transform 1 0 1360 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_12
timestamp 1714281807
transform 1 0 1288 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_13
timestamp 1714281807
transform 1 0 1264 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_14
timestamp 1714281807
transform 1 0 1360 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_15
timestamp 1714281807
transform 1 0 1472 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_16
timestamp 1714281807
transform 1 0 1416 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_17
timestamp 1714281807
transform 1 0 392 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_18
timestamp 1714281807
transform 1 0 392 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_19
timestamp 1714281807
transform 1 0 480 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_20
timestamp 1714281807
transform 1 0 464 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_21
timestamp 1714281807
transform 1 0 616 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_22
timestamp 1714281807
transform 1 0 704 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_23
timestamp 1714281807
transform 1 0 600 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_24
timestamp 1714281807
transform 1 0 496 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_25
timestamp 1714281807
transform 1 0 1880 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_26
timestamp 1714281807
transform 1 0 1624 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_27
timestamp 1714281807
transform 1 0 1688 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_28
timestamp 1714281807
transform 1 0 1960 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_29
timestamp 1714281807
transform 1 0 720 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_30
timestamp 1714281807
transform 1 0 664 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_31
timestamp 1714281807
transform 1 0 680 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_32
timestamp 1714281807
transform 1 0 728 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_33
timestamp 1714281807
transform 1 0 632 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_34
timestamp 1714281807
transform 1 0 968 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_35
timestamp 1714281807
transform 1 0 1040 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_36
timestamp 1714281807
transform 1 0 936 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_37
timestamp 1714281807
transform 1 0 1040 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_38
timestamp 1714281807
transform 1 0 824 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_39
timestamp 1714281807
transform 1 0 872 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_40
timestamp 1714281807
transform 1 0 736 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_41
timestamp 1714281807
transform 1 0 1904 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_42
timestamp 1714281807
transform 1 0 1768 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_43
timestamp 1714281807
transform 1 0 1560 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_44
timestamp 1714281807
transform 1 0 1272 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_45
timestamp 1714281807
transform 1 0 1176 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_46
timestamp 1714281807
transform 1 0 1208 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_47
timestamp 1714281807
transform 1 0 1208 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_48
timestamp 1714281807
transform 1 0 1248 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_49
timestamp 1714281807
transform 1 0 800 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_50
timestamp 1714281807
transform 1 0 672 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_51
timestamp 1714281807
transform 1 0 1400 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_52
timestamp 1714281807
transform 1 0 808 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_53
timestamp 1714281807
transform 1 0 496 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_54
timestamp 1714281807
transform 1 0 256 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_55
timestamp 1714281807
transform 1 0 248 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_56
timestamp 1714281807
transform 1 0 224 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_57
timestamp 1714281807
transform 1 0 256 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_58
timestamp 1714281807
transform 1 0 328 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_59
timestamp 1714281807
transform 1 0 496 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_60
timestamp 1714281807
transform 1 0 664 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_61
timestamp 1714281807
transform 1 0 640 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_62
timestamp 1714281807
transform 1 0 824 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_63
timestamp 1714281807
transform 1 0 568 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_64
timestamp 1714281807
transform 1 0 600 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_65
timestamp 1714281807
transform 1 0 560 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_66
timestamp 1714281807
transform 1 0 248 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_67
timestamp 1714281807
transform 1 0 696 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_68
timestamp 1714281807
transform 1 0 616 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_69
timestamp 1714281807
transform 1 0 632 0 1 570
box -8 -3 32 105
use NAND3X1  NAND3X1_0
timestamp 1714281807
transform 1 0 400 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_1
timestamp 1714281807
transform 1 0 2200 0 1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_2
timestamp 1714281807
transform 1 0 2744 0 -1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_3
timestamp 1714281807
transform 1 0 2424 0 1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_4
timestamp 1714281807
transform 1 0 2624 0 1 2570
box -8 -3 40 105
use NAND3X1  NAND3X1_5
timestamp 1714281807
transform 1 0 1568 0 -1 2770
box -8 -3 40 105
use NAND3X1  NAND3X1_6
timestamp 1714281807
transform 1 0 2176 0 -1 2770
box -8 -3 40 105
use NAND3X1  NAND3X1_7
timestamp 1714281807
transform 1 0 2024 0 1 2570
box -8 -3 40 105
use NAND3X1  NAND3X1_8
timestamp 1714281807
transform 1 0 2280 0 -1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_9
timestamp 1714281807
transform 1 0 2600 0 -1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_10
timestamp 1714281807
transform 1 0 1464 0 -1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_11
timestamp 1714281807
transform 1 0 1920 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_12
timestamp 1714281807
transform 1 0 1616 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_13
timestamp 1714281807
transform 1 0 2648 0 1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_14
timestamp 1714281807
transform 1 0 2368 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_15
timestamp 1714281807
transform 1 0 1688 0 1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_16
timestamp 1714281807
transform 1 0 1552 0 -1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_17
timestamp 1714281807
transform 1 0 1184 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_18
timestamp 1714281807
transform 1 0 1312 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_19
timestamp 1714281807
transform 1 0 928 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_20
timestamp 1714281807
transform 1 0 856 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_21
timestamp 1714281807
transform 1 0 664 0 1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_22
timestamp 1714281807
transform 1 0 1720 0 -1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_23
timestamp 1714281807
transform 1 0 1504 0 -1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_24
timestamp 1714281807
transform 1 0 1784 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_25
timestamp 1714281807
transform 1 0 624 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_26
timestamp 1714281807
transform 1 0 592 0 -1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_27
timestamp 1714281807
transform 1 0 536 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_28
timestamp 1714281807
transform 1 0 480 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_29
timestamp 1714281807
transform 1 0 640 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_30
timestamp 1714281807
transform 1 0 640 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_31
timestamp 1714281807
transform 1 0 952 0 -1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_32
timestamp 1714281807
transform 1 0 1000 0 -1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_33
timestamp 1714281807
transform 1 0 1184 0 1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_34
timestamp 1714281807
transform 1 0 1160 0 -1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_35
timestamp 1714281807
transform 1 0 1112 0 1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_36
timestamp 1714281807
transform 1 0 1048 0 -1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_37
timestamp 1714281807
transform 1 0 672 0 -1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_38
timestamp 1714281807
transform 1 0 1808 0 1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_39
timestamp 1714281807
transform 1 0 624 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_40
timestamp 1714281807
transform 1 0 552 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_41
timestamp 1714281807
transform 1 0 360 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_42
timestamp 1714281807
transform 1 0 320 0 -1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_43
timestamp 1714281807
transform 1 0 664 0 -1 170
box -8 -3 40 105
use NOR2X1  NOR2X1_0
timestamp 1714281807
transform 1 0 1064 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_1
timestamp 1714281807
transform 1 0 912 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_2
timestamp 1714281807
transform 1 0 776 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_3
timestamp 1714281807
transform 1 0 848 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_4
timestamp 1714281807
transform 1 0 456 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_5
timestamp 1714281807
transform 1 0 352 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_6
timestamp 1714281807
transform 1 0 352 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_7
timestamp 1714281807
transform 1 0 496 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_8
timestamp 1714281807
transform 1 0 952 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_9
timestamp 1714281807
transform 1 0 1008 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_10
timestamp 1714281807
transform 1 0 1168 0 1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_11
timestamp 1714281807
transform 1 0 1224 0 1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_12
timestamp 1714281807
transform 1 0 2472 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_13
timestamp 1714281807
transform 1 0 2432 0 1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_14
timestamp 1714281807
transform 1 0 2176 0 1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_15
timestamp 1714281807
transform 1 0 2288 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_16
timestamp 1714281807
transform 1 0 1768 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_17
timestamp 1714281807
transform 1 0 2376 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_18
timestamp 1714281807
transform 1 0 1624 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_19
timestamp 1714281807
transform 1 0 1640 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_20
timestamp 1714281807
transform 1 0 1376 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_21
timestamp 1714281807
transform 1 0 800 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_22
timestamp 1714281807
transform 1 0 872 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_23
timestamp 1714281807
transform 1 0 600 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_24
timestamp 1714281807
transform 1 0 816 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_25
timestamp 1714281807
transform 1 0 792 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_26
timestamp 1714281807
transform 1 0 1288 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_27
timestamp 1714281807
transform 1 0 2416 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_28
timestamp 1714281807
transform 1 0 2552 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_29
timestamp 1714281807
transform 1 0 2456 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_30
timestamp 1714281807
transform 1 0 2680 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_31
timestamp 1714281807
transform 1 0 2584 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_32
timestamp 1714281807
transform 1 0 2632 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_33
timestamp 1714281807
transform 1 0 2088 0 -1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_34
timestamp 1714281807
transform 1 0 2256 0 -1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_35
timestamp 1714281807
transform 1 0 2416 0 -1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_36
timestamp 1714281807
transform 1 0 1784 0 -1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_37
timestamp 1714281807
transform 1 0 1840 0 -1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_38
timestamp 1714281807
transform 1 0 2048 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_39
timestamp 1714281807
transform 1 0 2616 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_40
timestamp 1714281807
transform 1 0 2688 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_41
timestamp 1714281807
transform 1 0 2872 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_42
timestamp 1714281807
transform 1 0 1520 0 -1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_43
timestamp 1714281807
transform 1 0 1616 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_44
timestamp 1714281807
transform 1 0 1560 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_45
timestamp 1714281807
transform 1 0 2680 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_46
timestamp 1714281807
transform 1 0 2832 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_47
timestamp 1714281807
transform 1 0 2880 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_48
timestamp 1714281807
transform 1 0 2576 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_49
timestamp 1714281807
transform 1 0 2416 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_50
timestamp 1714281807
transform 1 0 2504 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_51
timestamp 1714281807
transform 1 0 2728 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_52
timestamp 1714281807
transform 1 0 2864 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_53
timestamp 1714281807
transform 1 0 2848 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_54
timestamp 1714281807
transform 1 0 2248 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_55
timestamp 1714281807
transform 1 0 2584 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_56
timestamp 1714281807
transform 1 0 2424 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_57
timestamp 1714281807
transform 1 0 1848 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_58
timestamp 1714281807
transform 1 0 2016 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_59
timestamp 1714281807
transform 1 0 2064 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_60
timestamp 1714281807
transform 1 0 1360 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_61
timestamp 1714281807
transform 1 0 1688 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_62
timestamp 1714281807
transform 1 0 1528 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_63
timestamp 1714281807
transform 1 0 1184 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_64
timestamp 1714281807
transform 1 0 992 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_65
timestamp 1714281807
transform 1 0 1032 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_66
timestamp 1714281807
transform 1 0 1088 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_67
timestamp 1714281807
transform 1 0 1072 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_68
timestamp 1714281807
transform 1 0 1040 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_69
timestamp 1714281807
transform 1 0 1792 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_70
timestamp 1714281807
transform 1 0 1672 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_71
timestamp 1714281807
transform 1 0 1768 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_72
timestamp 1714281807
transform 1 0 1736 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_73
timestamp 1714281807
transform 1 0 1536 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_74
timestamp 1714281807
transform 1 0 1576 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_75
timestamp 1714281807
transform 1 0 2088 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_76
timestamp 1714281807
transform 1 0 2032 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_77
timestamp 1714281807
transform 1 0 2264 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_78
timestamp 1714281807
transform 1 0 2808 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_79
timestamp 1714281807
transform 1 0 2816 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_80
timestamp 1714281807
transform 1 0 2824 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_81
timestamp 1714281807
transform 1 0 2112 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_82
timestamp 1714281807
transform 1 0 2264 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_83
timestamp 1714281807
transform 1 0 2392 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_84
timestamp 1714281807
transform 1 0 1736 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_85
timestamp 1714281807
transform 1 0 1952 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_86
timestamp 1714281807
transform 1 0 2016 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_87
timestamp 1714281807
transform 1 0 2520 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_88
timestamp 1714281807
transform 1 0 2768 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_89
timestamp 1714281807
transform 1 0 2808 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_90
timestamp 1714281807
transform 1 0 1568 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_91
timestamp 1714281807
transform 1 0 1624 0 -1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_92
timestamp 1714281807
transform 1 0 1560 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_93
timestamp 1714281807
transform 1 0 2504 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_94
timestamp 1714281807
transform 1 0 2816 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_95
timestamp 1714281807
transform 1 0 2712 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_96
timestamp 1714281807
transform 1 0 2232 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_97
timestamp 1714281807
transform 1 0 2480 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_98
timestamp 1714281807
transform 1 0 2408 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_99
timestamp 1714281807
transform 1 0 2720 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_100
timestamp 1714281807
transform 1 0 2816 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_101
timestamp 1714281807
transform 1 0 2792 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_102
timestamp 1714281807
transform 1 0 2304 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_103
timestamp 1714281807
transform 1 0 2520 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_104
timestamp 1714281807
transform 1 0 2552 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_105
timestamp 1714281807
transform 1 0 1840 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_106
timestamp 1714281807
transform 1 0 2200 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_107
timestamp 1714281807
transform 1 0 2104 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_108
timestamp 1714281807
transform 1 0 1952 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_109
timestamp 1714281807
transform 1 0 2032 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_110
timestamp 1714281807
transform 1 0 1672 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_111
timestamp 1714281807
transform 1 0 1464 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_112
timestamp 1714281807
transform 1 0 1632 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_113
timestamp 1714281807
transform 1 0 1472 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_114
timestamp 1714281807
transform 1 0 1544 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_115
timestamp 1714281807
transform 1 0 1432 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_116
timestamp 1714281807
transform 1 0 1472 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_117
timestamp 1714281807
transform 1 0 2104 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_118
timestamp 1714281807
transform 1 0 2032 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_119
timestamp 1714281807
transform 1 0 1992 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_120
timestamp 1714281807
transform 1 0 1880 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_121
timestamp 1714281807
transform 1 0 2112 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_122
timestamp 1714281807
transform 1 0 2088 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_123
timestamp 1714281807
transform 1 0 984 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_124
timestamp 1714281807
transform 1 0 480 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_125
timestamp 1714281807
transform 1 0 504 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_126
timestamp 1714281807
transform 1 0 216 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_127
timestamp 1714281807
transform 1 0 888 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_128
timestamp 1714281807
transform 1 0 280 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_129
timestamp 1714281807
transform 1 0 256 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_130
timestamp 1714281807
transform 1 0 736 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_131
timestamp 1714281807
transform 1 0 792 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_132
timestamp 1714281807
transform 1 0 496 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_133
timestamp 1714281807
transform 1 0 680 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_134
timestamp 1714281807
transform 1 0 568 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_135
timestamp 1714281807
transform 1 0 400 0 -1 770
box -8 -3 32 105
use OAI21X1  OAI21X1_0
timestamp 1714281807
transform 1 0 808 0 -1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_1
timestamp 1714281807
transform 1 0 648 0 -1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_2
timestamp 1714281807
transform 1 0 264 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_3
timestamp 1714281807
transform 1 0 440 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_4
timestamp 1714281807
transform 1 0 648 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_5
timestamp 1714281807
transform 1 0 808 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_6
timestamp 1714281807
transform 1 0 2488 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_7
timestamp 1714281807
transform 1 0 2568 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_8
timestamp 1714281807
transform 1 0 2288 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_9
timestamp 1714281807
transform 1 0 2096 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_10
timestamp 1714281807
transform 1 0 2040 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_11
timestamp 1714281807
transform 1 0 1856 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_12
timestamp 1714281807
transform 1 0 1496 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_13
timestamp 1714281807
transform 1 0 1680 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_14
timestamp 1714281807
transform 1 0 1408 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_15
timestamp 1714281807
transform 1 0 1048 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_16
timestamp 1714281807
transform 1 0 1096 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_17
timestamp 1714281807
transform 1 0 1264 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_18
timestamp 1714281807
transform 1 0 1104 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_19
timestamp 1714281807
transform 1 0 1088 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_20
timestamp 1714281807
transform 1 0 1152 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_21
timestamp 1714281807
transform 1 0 1824 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_22
timestamp 1714281807
transform 1 0 1608 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_23
timestamp 1714281807
transform 1 0 1832 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_24
timestamp 1714281807
transform 1 0 1552 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_25
timestamp 1714281807
transform 1 0 1560 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_26
timestamp 1714281807
transform 1 0 1736 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_27
timestamp 1714281807
transform 1 0 2368 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_28
timestamp 1714281807
transform 1 0 2416 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_29
timestamp 1714281807
transform 1 0 2408 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_30
timestamp 1714281807
transform 1 0 2840 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_31
timestamp 1714281807
transform 1 0 2752 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_32
timestamp 1714281807
transform 1 0 2880 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_33
timestamp 1714281807
transform 1 0 2288 0 -1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_34
timestamp 1714281807
transform 1 0 2056 0 -1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_35
timestamp 1714281807
transform 1 0 2416 0 -1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_36
timestamp 1714281807
transform 1 0 1872 0 -1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_37
timestamp 1714281807
transform 1 0 1760 0 -1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_38
timestamp 1714281807
transform 1 0 1960 0 -1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_39
timestamp 1714281807
transform 1 0 2720 0 -1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_40
timestamp 1714281807
transform 1 0 2504 0 -1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_41
timestamp 1714281807
transform 1 0 2800 0 -1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_42
timestamp 1714281807
transform 1 0 1296 0 1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_43
timestamp 1714281807
transform 1 0 1440 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_44
timestamp 1714281807
transform 1 0 1360 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_45
timestamp 1714281807
transform 1 0 2824 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_46
timestamp 1714281807
transform 1 0 2624 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_47
timestamp 1714281807
transform 1 0 2832 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_48
timestamp 1714281807
transform 1 0 2336 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_49
timestamp 1714281807
transform 1 0 2136 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_50
timestamp 1714281807
transform 1 0 2312 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_51
timestamp 1714281807
transform 1 0 2824 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_52
timestamp 1714281807
transform 1 0 2736 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_53
timestamp 1714281807
transform 1 0 2832 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_54
timestamp 1714281807
transform 1 0 920 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_55
timestamp 1714281807
transform 1 0 904 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_56
timestamp 1714281807
transform 1 0 936 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_57
timestamp 1714281807
transform 1 0 1008 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_58
timestamp 1714281807
transform 1 0 504 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_59
timestamp 1714281807
transform 1 0 576 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_60
timestamp 1714281807
transform 1 0 528 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_61
timestamp 1714281807
transform 1 0 336 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_62
timestamp 1714281807
transform 1 0 2416 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_63
timestamp 1714281807
transform 1 0 2440 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_64
timestamp 1714281807
transform 1 0 2288 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_65
timestamp 1714281807
transform 1 0 2400 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_66
timestamp 1714281807
transform 1 0 2472 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_67
timestamp 1714281807
transform 1 0 2312 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_68
timestamp 1714281807
transform 1 0 2016 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_69
timestamp 1714281807
transform 1 0 2088 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_70
timestamp 1714281807
transform 1 0 1776 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_71
timestamp 1714281807
transform 1 0 1752 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_72
timestamp 1714281807
transform 1 0 1960 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_73
timestamp 1714281807
transform 1 0 1856 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_74
timestamp 1714281807
transform 1 0 1400 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_75
timestamp 1714281807
transform 1 0 1672 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_76
timestamp 1714281807
transform 1 0 1400 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_77
timestamp 1714281807
transform 1 0 1416 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_78
timestamp 1714281807
transform 1 0 1544 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_79
timestamp 1714281807
transform 1 0 1496 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_80
timestamp 1714281807
transform 1 0 1440 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_81
timestamp 1714281807
transform 1 0 1376 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_82
timestamp 1714281807
transform 1 0 1528 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_83
timestamp 1714281807
transform 1 0 1984 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_84
timestamp 1714281807
transform 1 0 1960 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_85
timestamp 1714281807
transform 1 0 2000 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_86
timestamp 1714281807
transform 1 0 2136 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_87
timestamp 1714281807
transform 1 0 2080 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_88
timestamp 1714281807
transform 1 0 1976 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_89
timestamp 1714281807
transform 1 0 2688 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_90
timestamp 1714281807
transform 1 0 2592 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_91
timestamp 1714281807
transform 1 0 2464 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_92
timestamp 1714281807
transform 1 0 2608 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_93
timestamp 1714281807
transform 1 0 2640 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_94
timestamp 1714281807
transform 1 0 2488 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_95
timestamp 1714281807
transform 1 0 1952 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_96
timestamp 1714281807
transform 1 0 1872 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_97
timestamp 1714281807
transform 1 0 1776 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_98
timestamp 1714281807
transform 1 0 1624 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_99
timestamp 1714281807
transform 1 0 2328 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_100
timestamp 1714281807
transform 1 0 2200 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_101
timestamp 1714281807
transform 1 0 2112 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_102
timestamp 1714281807
transform 1 0 2736 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_103
timestamp 1714281807
transform 1 0 2744 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_104
timestamp 1714281807
transform 1 0 2672 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_105
timestamp 1714281807
transform 1 0 2344 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_106
timestamp 1714281807
transform 1 0 2136 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_107
timestamp 1714281807
transform 1 0 2128 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_108
timestamp 1714281807
transform 1 0 576 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_109
timestamp 1714281807
transform 1 0 432 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_110
timestamp 1714281807
transform 1 0 392 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_111
timestamp 1714281807
transform 1 0 240 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_112
timestamp 1714281807
transform 1 0 264 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_113
timestamp 1714281807
transform 1 0 312 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_114
timestamp 1714281807
transform 1 0 744 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_115
timestamp 1714281807
transform 1 0 392 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_116
timestamp 1714281807
transform 1 0 712 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_117
timestamp 1714281807
transform 1 0 544 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_118
timestamp 1714281807
transform 1 0 648 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_119
timestamp 1714281807
transform 1 0 856 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_120
timestamp 1714281807
transform 1 0 1256 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_121
timestamp 1714281807
transform 1 0 896 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_122
timestamp 1714281807
transform 1 0 720 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_123
timestamp 1714281807
transform 1 0 896 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_124
timestamp 1714281807
transform 1 0 824 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_125
timestamp 1714281807
transform 1 0 984 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_126
timestamp 1714281807
transform 1 0 1280 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_127
timestamp 1714281807
transform 1 0 1136 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_128
timestamp 1714281807
transform 1 0 1160 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_129
timestamp 1714281807
transform 1 0 1128 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_130
timestamp 1714281807
transform 1 0 2728 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_131
timestamp 1714281807
transform 1 0 2720 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_132
timestamp 1714281807
transform 1 0 2704 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_133
timestamp 1714281807
transform 1 0 1832 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_134
timestamp 1714281807
transform 1 0 680 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_135
timestamp 1714281807
transform 1 0 752 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_136
timestamp 1714281807
transform 1 0 472 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_137
timestamp 1714281807
transform 1 0 488 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_138
timestamp 1714281807
transform 1 0 392 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_139
timestamp 1714281807
transform 1 0 496 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_140
timestamp 1714281807
transform 1 0 416 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_141
timestamp 1714281807
transform 1 0 728 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_142
timestamp 1714281807
transform 1 0 864 0 -1 170
box -8 -3 34 105
use OAI22X1  OAI22X1_0
timestamp 1714281807
transform 1 0 848 0 1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_1
timestamp 1714281807
transform 1 0 944 0 -1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_2
timestamp 1714281807
transform 1 0 1104 0 -1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_3
timestamp 1714281807
transform 1 0 1144 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_4
timestamp 1714281807
transform 1 0 1072 0 1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_5
timestamp 1714281807
transform 1 0 760 0 1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_6
timestamp 1714281807
transform 1 0 592 0 -1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_7
timestamp 1714281807
transform 1 0 536 0 1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_8
timestamp 1714281807
transform 1 0 528 0 -1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_9
timestamp 1714281807
transform 1 0 368 0 -1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_10
timestamp 1714281807
transform 1 0 504 0 -1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_11
timestamp 1714281807
transform 1 0 256 0 1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_12
timestamp 1714281807
transform 1 0 272 0 -1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_13
timestamp 1714281807
transform 1 0 424 0 1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_14
timestamp 1714281807
transform 1 0 200 0 -1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_15
timestamp 1714281807
transform 1 0 248 0 1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_16
timestamp 1714281807
transform 1 0 1064 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_17
timestamp 1714281807
transform 1 0 944 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_18
timestamp 1714281807
transform 1 0 1440 0 1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_19
timestamp 1714281807
transform 1 0 856 0 -1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_20
timestamp 1714281807
transform 1 0 848 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_21
timestamp 1714281807
transform 1 0 1088 0 -1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_22
timestamp 1714281807
transform 1 0 416 0 1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_23
timestamp 1714281807
transform 1 0 408 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_24
timestamp 1714281807
transform 1 0 256 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_25
timestamp 1714281807
transform 1 0 432 0 1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_26
timestamp 1714281807
transform 1 0 504 0 1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_27
timestamp 1714281807
transform 1 0 584 0 1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_28
timestamp 1714281807
transform 1 0 672 0 1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_29
timestamp 1714281807
transform 1 0 520 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_30
timestamp 1714281807
transform 1 0 528 0 -1 1170
box -8 -3 46 105
use OAI22X1  OAI22X1_31
timestamp 1714281807
transform 1 0 480 0 -1 370
box -8 -3 46 105
use OR2X1  OR2X1_0
timestamp 1714281807
transform 1 0 864 0 1 970
box -8 -3 40 105
use OR2X1  OR2X1_1
timestamp 1714281807
transform 1 0 944 0 -1 1170
box -8 -3 40 105
use OR2X1  OR2X1_2
timestamp 1714281807
transform 1 0 936 0 1 1170
box -8 -3 40 105
use OR2X1  OR2X1_3
timestamp 1714281807
transform 1 0 1984 0 1 1370
box -8 -3 40 105
use OR2X1  OR2X1_4
timestamp 1714281807
transform 1 0 960 0 -1 2370
box -8 -3 40 105
use OR2X1  OR2X1_5
timestamp 1714281807
transform 1 0 728 0 -1 770
box -8 -3 40 105
use OR2X1  OR2X1_6
timestamp 1714281807
transform 1 0 336 0 -1 770
box -8 -3 40 105
use OR2X2  OR2X2_0
timestamp 1714281807
transform 1 0 704 0 1 2370
box -7 -3 35 105
use top_module_VIA0  top_module_VIA0_0
timestamp 1714281807
transform 1 0 3056 0 1 3017
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_1
timestamp 1714281807
transform 1 0 3056 0 1 23
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_2
timestamp 1714281807
transform 1 0 24 0 1 3017
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_3
timestamp 1714281807
transform 1 0 24 0 1 23
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_4
timestamp 1714281807
transform 1 0 3032 0 1 2993
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_5
timestamp 1714281807
transform 1 0 3032 0 1 47
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_6
timestamp 1714281807
transform 1 0 48 0 1 2993
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_7
timestamp 1714281807
transform 1 0 48 0 1 47
box -10 -10 10 10
use top_module_VIA1  top_module_VIA1_0
timestamp 1714281807
transform 1 0 3056 0 1 2870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_1
timestamp 1714281807
transform 1 0 3056 0 1 2670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_2
timestamp 1714281807
transform 1 0 3056 0 1 2470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_3
timestamp 1714281807
transform 1 0 3056 0 1 2270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_4
timestamp 1714281807
transform 1 0 3056 0 1 2070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_5
timestamp 1714281807
transform 1 0 3056 0 1 1870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_6
timestamp 1714281807
transform 1 0 3056 0 1 1670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_7
timestamp 1714281807
transform 1 0 3056 0 1 1470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_8
timestamp 1714281807
transform 1 0 3056 0 1 1270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_9
timestamp 1714281807
transform 1 0 3056 0 1 1070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_10
timestamp 1714281807
transform 1 0 3056 0 1 870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_11
timestamp 1714281807
transform 1 0 3056 0 1 670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_12
timestamp 1714281807
transform 1 0 3056 0 1 470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_13
timestamp 1714281807
transform 1 0 3056 0 1 270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_14
timestamp 1714281807
transform 1 0 3056 0 1 70
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_15
timestamp 1714281807
transform 1 0 24 0 1 2870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_16
timestamp 1714281807
transform 1 0 24 0 1 2670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_17
timestamp 1714281807
transform 1 0 24 0 1 2470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_18
timestamp 1714281807
transform 1 0 24 0 1 2270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_19
timestamp 1714281807
transform 1 0 24 0 1 2070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_20
timestamp 1714281807
transform 1 0 24 0 1 1870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_21
timestamp 1714281807
transform 1 0 24 0 1 1670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_22
timestamp 1714281807
transform 1 0 24 0 1 1470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_23
timestamp 1714281807
transform 1 0 24 0 1 1270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_24
timestamp 1714281807
transform 1 0 24 0 1 1070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_25
timestamp 1714281807
transform 1 0 24 0 1 870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_26
timestamp 1714281807
transform 1 0 24 0 1 670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_27
timestamp 1714281807
transform 1 0 24 0 1 470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_28
timestamp 1714281807
transform 1 0 24 0 1 270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_29
timestamp 1714281807
transform 1 0 24 0 1 70
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_30
timestamp 1714281807
transform 1 0 48 0 1 170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_31
timestamp 1714281807
transform 1 0 48 0 1 370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_32
timestamp 1714281807
transform 1 0 48 0 1 570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_33
timestamp 1714281807
transform 1 0 48 0 1 770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_34
timestamp 1714281807
transform 1 0 48 0 1 970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_35
timestamp 1714281807
transform 1 0 48 0 1 1170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_36
timestamp 1714281807
transform 1 0 48 0 1 1370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_37
timestamp 1714281807
transform 1 0 48 0 1 1570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_38
timestamp 1714281807
transform 1 0 48 0 1 1770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_39
timestamp 1714281807
transform 1 0 48 0 1 1970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_40
timestamp 1714281807
transform 1 0 48 0 1 2170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_41
timestamp 1714281807
transform 1 0 48 0 1 2370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_42
timestamp 1714281807
transform 1 0 48 0 1 2570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_43
timestamp 1714281807
transform 1 0 48 0 1 2770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_44
timestamp 1714281807
transform 1 0 48 0 1 2970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_45
timestamp 1714281807
transform 1 0 3032 0 1 170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_46
timestamp 1714281807
transform 1 0 3032 0 1 370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_47
timestamp 1714281807
transform 1 0 3032 0 1 570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_48
timestamp 1714281807
transform 1 0 3032 0 1 770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_49
timestamp 1714281807
transform 1 0 3032 0 1 970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_50
timestamp 1714281807
transform 1 0 3032 0 1 1170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_51
timestamp 1714281807
transform 1 0 3032 0 1 1370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_52
timestamp 1714281807
transform 1 0 3032 0 1 1570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_53
timestamp 1714281807
transform 1 0 3032 0 1 1770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_54
timestamp 1714281807
transform 1 0 3032 0 1 1970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_55
timestamp 1714281807
transform 1 0 3032 0 1 2170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_56
timestamp 1714281807
transform 1 0 3032 0 1 2370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_57
timestamp 1714281807
transform 1 0 3032 0 1 2570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_58
timestamp 1714281807
transform 1 0 3032 0 1 2770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_59
timestamp 1714281807
transform 1 0 3032 0 1 2970
box -10 -3 10 3
use XNOR2X1  XNOR2X1_0
timestamp 1714281807
transform 1 0 680 0 1 2770
box -8 -3 64 105
use XNOR2X1  XNOR2X1_1
timestamp 1714281807
transform 1 0 896 0 -1 2970
box -8 -3 64 105
use XNOR2X1  XNOR2X1_2
timestamp 1714281807
transform 1 0 1944 0 1 2170
box -8 -3 64 105
use XNOR2X1  XNOR2X1_3
timestamp 1714281807
transform 1 0 1864 0 1 2170
box -8 -3 64 105
use XNOR2X1  XNOR2X1_4
timestamp 1714281807
transform 1 0 1816 0 -1 1970
box -8 -3 64 105
use XOR2X1  XOR2X1_0
timestamp 1714281807
transform 1 0 864 0 1 2770
box -8 -3 64 105
use XOR2X1  XOR2X1_1
timestamp 1714281807
transform 1 0 2672 0 -1 1370
box -8 -3 64 105
use XOR2X1  XOR2X1_2
timestamp 1714281807
transform 1 0 2792 0 -1 1370
box -8 -3 64 105
use XOR2X1  XOR2X1_3
timestamp 1714281807
transform 1 0 2848 0 -1 1370
box -8 -3 64 105
use XOR2X1  XOR2X1_4
timestamp 1714281807
transform 1 0 2432 0 -1 1170
box -8 -3 64 105
use XOR2X1  XOR2X1_5
timestamp 1714281807
transform 1 0 2360 0 1 1170
box -8 -3 64 105
use XOR2X1  XOR2X1_6
timestamp 1714281807
transform 1 0 2376 0 -1 1170
box -8 -3 64 105
use XOR2X1  XOR2X1_7
timestamp 1714281807
transform 1 0 2568 0 -1 2770
box -8 -3 64 105
use XOR2X1  XOR2X1_8
timestamp 1714281807
transform 1 0 2632 0 -1 2770
box -8 -3 64 105
use XOR2X1  XOR2X1_9
timestamp 1714281807
transform 1 0 2848 0 1 2570
box -8 -3 64 105
use XOR2X1  XOR2X1_10
timestamp 1714281807
transform 1 0 1496 0 1 2770
box -8 -3 64 105
use XOR2X1  XOR2X1_11
timestamp 1714281807
transform 1 0 1576 0 1 2570
box -8 -3 64 105
use XOR2X1  XOR2X1_12
timestamp 1714281807
transform 1 0 1504 0 -1 2770
box -8 -3 64 105
use XOR2X1  XOR2X1_13
timestamp 1714281807
transform 1 0 2096 0 -1 2770
box -8 -3 64 105
use XOR2X1  XOR2X1_14
timestamp 1714281807
transform 1 0 2216 0 -1 2770
box -8 -3 64 105
use XOR2X1  XOR2X1_15
timestamp 1714281807
transform 1 0 2344 0 -1 2770
box -8 -3 64 105
use XOR2X1  XOR2X1_16
timestamp 1714281807
transform 1 0 1800 0 -1 2770
box -8 -3 64 105
use XOR2X1  XOR2X1_17
timestamp 1714281807
transform 1 0 1856 0 1 2570
box -8 -3 64 105
use XOR2X1  XOR2X1_18
timestamp 1714281807
transform 1 0 1968 0 1 2570
box -8 -3 64 105
use XOR2X1  XOR2X1_19
timestamp 1714281807
transform 1 0 2328 0 -1 2170
box -8 -3 64 105
use XOR2X1  XOR2X1_20
timestamp 1714281807
transform 1 0 2304 0 -1 1970
box -8 -3 64 105
use XOR2X1  XOR2X1_21
timestamp 1714281807
transform 1 0 2240 0 -1 1770
box -8 -3 64 105
use XOR2X1  XOR2X1_22
timestamp 1714281807
transform 1 0 2672 0 1 2170
box -8 -3 64 105
use XOR2X1  XOR2X1_23
timestamp 1714281807
transform 1 0 2624 0 1 1970
box -8 -3 64 105
use XOR2X1  XOR2X1_24
timestamp 1714281807
transform 1 0 2632 0 -1 2170
box -8 -3 64 105
use XOR2X1  XOR2X1_25
timestamp 1714281807
transform 1 0 2216 0 -1 370
box -8 -3 64 105
use XOR2X1  XOR2X1_26
timestamp 1714281807
transform 1 0 1728 0 -1 370
box -8 -3 64 105
use XOR2X1  XOR2X1_27
timestamp 1714281807
transform 1 0 1968 0 -1 370
box -8 -3 64 105
use XOR2X1  XOR2X1_28
timestamp 1714281807
transform 1 0 1784 0 -1 370
box -8 -3 64 105
use XOR2X1  XOR2X1_29
timestamp 1714281807
transform 1 0 1320 0 -1 370
box -8 -3 64 105
use XOR2X1  XOR2X1_30
timestamp 1714281807
transform 1 0 1536 0 -1 370
box -8 -3 64 105
use XOR2X1  XOR2X1_31
timestamp 1714281807
transform 1 0 2872 0 1 370
box -8 -3 64 105
use XOR2X1  XOR2X1_32
timestamp 1714281807
transform 1 0 2592 0 1 370
box -8 -3 64 105
use XOR2X1  XOR2X1_33
timestamp 1714281807
transform 1 0 2656 0 -1 570
box -8 -3 64 105
use XOR2X1  XOR2X1_34
timestamp 1714281807
transform 1 0 2640 0 -1 370
box -8 -3 64 105
use XOR2X1  XOR2X1_35
timestamp 1714281807
transform 1 0 2152 0 -1 370
box -8 -3 64 105
use XOR2X1  XOR2X1_36
timestamp 1714281807
transform 1 0 2408 0 -1 370
box -8 -3 64 105
use XOR2X1  XOR2X1_37
timestamp 1714281807
transform 1 0 1352 0 -1 1170
box -8 -3 64 105
use XOR2X1  XOR2X1_38
timestamp 1714281807
transform 1 0 1672 0 1 1370
box -8 -3 64 105
use XOR2X1  XOR2X1_39
timestamp 1714281807
transform 1 0 1760 0 -1 1170
box -8 -3 64 105
use XOR2X1  XOR2X1_40
timestamp 1714281807
transform 1 0 1672 0 -1 1370
box -8 -3 64 105
use XOR2X1  XOR2X1_41
timestamp 1714281807
transform 1 0 1800 0 1 1570
box -8 -3 64 105
use XOR2X1  XOR2X1_42
timestamp 1714281807
transform 1 0 1608 0 1 1570
box -8 -3 64 105
use XOR2X1  XOR2X1_43
timestamp 1714281807
transform 1 0 1328 0 1 370
box -8 -3 64 105
use XOR2X1  XOR2X1_44
timestamp 1714281807
transform 1 0 1112 0 1 570
box -8 -3 64 105
use XOR2X1  XOR2X1_45
timestamp 1714281807
transform 1 0 1128 0 -1 570
box -8 -3 64 105
use XOR2X1  XOR2X1_46
timestamp 1714281807
transform 1 0 1200 0 -1 570
box -8 -3 64 105
use XOR2X1  XOR2X1_47
timestamp 1714281807
transform 1 0 1592 0 -1 970
box -8 -3 64 105
use XOR2X1  XOR2X1_48
timestamp 1714281807
transform 1 0 1240 0 1 770
box -8 -3 64 105
use XOR2X1  XOR2X1_49
timestamp 1714281807
transform 1 0 1504 0 1 2170
box -8 -3 64 105
use XOR2X1  XOR2X1_50
timestamp 1714281807
transform 1 0 1568 0 1 1970
box -8 -3 64 105
use XOR2X1  XOR2X1_51
timestamp 1714281807
transform 1 0 568 0 1 370
box -8 -3 64 105
<< labels >>
rlabel metal2 1588 3038 1588 3038 4 in_clka
rlabel metal2 1572 1 1572 1 4 in_clkb
rlabel metal3 2 2195 2 2195 4 in_restart
rlabel metal3 2 1455 2 1455 4 in_new_game
rlabel metal2 340 1 340 1 4 in_enter
rlabel metal3 2 1135 2 1135 4 in_diff_cell_val[1]
rlabel metal3 2 1075 2 1075 4 in_diff_cell_val[0]
rlabel metal2 884 1 884 1 4 out_solved
rlabel metal2 508 1 508 1 4 out_state[3]
rlabel metal2 476 1 476 1 4 out_state[2]
rlabel metal2 492 1 492 1 4 out_state[1]
rlabel metal2 652 1 652 1 4 out_state[0]
rlabel metal2 1508 3038 1508 3038 4 in_rand_setup[3]
rlabel metal2 1748 3038 1748 3038 4 in_rand_setup[2]
rlabel metal2 1628 3038 1628 3038 4 in_rand_setup[1]
rlabel metal2 1572 3038 1572 3038 4 in_rand_setup[0]
rlabel metal3 2 2065 2 2065 4 in_rand_A[3]
rlabel metal3 2 1775 2 1775 4 in_rand_A[2]
rlabel metal3 2 2105 2 2105 4 in_rand_A[1]
rlabel metal3 2 2125 2 2125 4 in_rand_A[0]
rlabel metal2 1132 3038 1132 3038 4 in_rand_B[3]
rlabel metal2 1116 3038 1116 3038 4 in_rand_B[2]
rlabel metal2 908 3038 908 3038 4 in_rand_B[1]
rlabel metal2 1020 3038 1020 3038 4 in_rand_B[0]
rlabel metal3 2 855 2 855 4 out_gen_rand_flag
rlabel metal3 2 875 2 875 4 out_set_board_flag
rlabel metal3 2 975 2 975 4 out_set_diff_flag
rlabel metal3 2 895 2 895 4 out_row_flag
rlabel metal3 2 915 2 915 4 out_col_flag
rlabel metal2 868 1 868 1 4 out_val_flag
rlabel metal2 932 1 932 1 4 out_check_flag
rlabel metal2 1468 3038 1468 3038 4 out_fill_flag[15]
rlabel metal2 1484 3038 1484 3038 4 out_fill_flag[14]
rlabel metal2 1548 3038 1548 3038 4 out_fill_flag[13]
rlabel metal2 1452 3038 1452 3038 4 out_fill_flag[12]
rlabel metal2 828 3038 828 3038 4 out_fill_flag[11]
rlabel metal2 804 3038 804 3038 4 out_fill_flag[10]
rlabel metal2 1524 3038 1524 3038 4 out_fill_flag[9]
rlabel metal3 2 1725 2 1725 4 out_fill_flag[8]
rlabel metal3 2 1815 2 1815 4 out_fill_flag[7]
rlabel metal3 2 1525 2 1525 4 out_fill_flag[6]
rlabel metal3 2 1325 2 1325 4 out_fill_flag[5]
rlabel metal3 2 1015 2 1015 4 out_fill_flag[4]
rlabel metal3 2 2015 2 2015 4 out_fill_flag[3]
rlabel metal3 2 2145 2 2145 4 out_fill_flag[2]
rlabel metal3 2 2215 2 2215 4 out_fill_flag[1]
rlabel metal3 2 815 2 815 4 out_fill_flag[0]
rlabel metal2 1804 3038 1804 3038 4 out_user_board_0[2]
rlabel metal2 1668 1 1668 1 4 out_user_board_0[1]
rlabel metal2 1676 3038 1676 3038 4 out_user_board_0[0]
rlabel metal3 3077 1565 3077 1565 4 out_user_board_1[2]
rlabel metal2 1716 1 1716 1 4 out_user_board_1[1]
rlabel metal2 1820 1 1820 1 4 out_user_board_1[0]
rlabel metal2 1156 1 1156 1 4 out_user_board_2[2]
rlabel metal2 996 1 996 1 4 out_user_board_2[1]
rlabel metal2 1012 1 1012 1 4 out_user_board_2[0]
rlabel metal2 1140 1 1140 1 4 out_user_board_3[2]
rlabel metal2 1036 1 1036 1 4 out_user_board_3[1]
rlabel metal2 980 1 980 1 4 out_user_board_3[0]
rlabel metal2 1332 1 1332 1 4 out_user_board_4[2]
rlabel metal2 1684 1 1684 1 4 out_user_board_4[1]
rlabel metal2 1508 1 1508 1 4 out_user_board_4[0]
rlabel metal2 1836 1 1836 1 4 out_user_board_5[2]
rlabel metal2 1980 1 1980 1 4 out_user_board_5[1]
rlabel metal2 2220 1 2220 1 4 out_user_board_5[0]
rlabel metal2 2388 1 2388 1 4 out_user_board_6[2]
rlabel metal2 2708 1 2708 1 4 out_user_board_6[1]
rlabel metal2 2564 1 2564 1 4 out_user_board_6[0]
rlabel metal2 2844 1 2844 1 4 out_user_board_7[2]
rlabel metal3 3077 125 3077 125 4 out_user_board_7[1]
rlabel metal3 3077 215 3077 215 4 out_user_board_7[0]
rlabel metal3 3077 1015 3077 1015 4 out_user_board_8[2]
rlabel metal3 3077 995 3077 995 4 out_user_board_8[1]
rlabel metal3 3077 1105 3077 1105 4 out_user_board_8[0]
rlabel metal3 3077 1145 3077 1145 4 out_user_board_9[2]
rlabel metal3 3077 1085 3077 1085 4 out_user_board_9[1]
rlabel metal3 3077 1035 3077 1035 4 out_user_board_9[0]
rlabel metal2 1660 3038 1660 3038 4 out_user_board_10[2]
rlabel metal2 1764 3038 1764 3038 4 out_user_board_10[1]
rlabel metal2 1644 3038 1644 3038 4 out_user_board_10[0]
rlabel metal2 2660 3038 2660 3038 4 out_user_board_11[2]
rlabel metal2 2764 3038 2764 3038 4 out_user_board_11[1]
rlabel metal2 2868 3038 2868 3038 4 out_user_board_11[0]
rlabel metal2 1780 3038 1780 3038 4 out_user_board_12[2]
rlabel metal2 1972 3038 1972 3038 4 out_user_board_12[1]
rlabel metal2 2052 3038 2052 3038 4 out_user_board_12[0]
rlabel metal2 2220 3038 2220 3038 4 out_user_board_13[2]
rlabel metal2 2388 3038 2388 3038 4 out_user_board_13[1]
rlabel metal2 2556 3038 2556 3038 4 out_user_board_13[0]
rlabel metal3 3077 2345 3077 2345 4 out_user_board_14[2]
rlabel metal3 3077 2015 3077 2015 4 out_user_board_14[1]
rlabel metal3 3077 2215 3077 2215 4 out_user_board_14[0]
rlabel metal3 3077 2105 3077 2105 4 out_user_board_15[2]
rlabel metal3 3077 1835 3077 1835 4 out_user_board_15[1]
rlabel metal3 3077 1705 3077 1705 4 out_user_board_15[0]
rlabel metal3 3077 1525 3077 1525 4 out_real_board_0[2]
rlabel metal3 3077 1415 3077 1415 4 out_real_board_0[1]
rlabel metal3 3077 1505 3077 1505 4 out_real_board_0[0]
rlabel metal3 3077 1215 3077 1215 4 out_real_board_1[2]
rlabel metal3 3077 925 3077 925 4 out_real_board_1[1]
rlabel metal3 3077 1125 3077 1125 4 out_real_board_1[0]
rlabel metal2 1604 1 1604 1 4 out_real_board_2[2]
rlabel metal2 1556 1 1556 1 4 out_real_board_2[1]
rlabel metal2 1620 1 1620 1 4 out_real_board_2[0]
rlabel metal2 1588 1 1588 1 4 out_real_board_3[2]
rlabel metal2 1748 1 1748 1 4 out_real_board_3[1]
rlabel metal2 1636 1 1636 1 4 out_real_board_3[0]
rlabel metal2 2100 1 2100 1 4 out_real_board_4[2]
rlabel metal2 2164 1 2164 1 4 out_real_board_4[1]
rlabel metal2 1652 1 1652 1 4 out_real_board_4[0]
rlabel metal2 1916 1 1916 1 4 out_real_board_5[2]
rlabel metal2 2252 1 2252 1 4 out_real_board_5[1]
rlabel metal2 2268 1 2268 1 4 out_real_board_5[0]
rlabel metal3 3077 725 3077 725 4 out_real_board_6[2]
rlabel metal3 3077 705 3077 705 4 out_real_board_6[1]
rlabel metal3 3077 615 3077 615 4 out_real_board_6[0]
rlabel metal3 3077 595 3077 595 4 out_real_board_7[2]
rlabel metal3 3077 815 3077 815 4 out_real_board_7[1]
rlabel metal3 3077 905 3077 905 4 out_real_board_7[0]
rlabel metal2 2204 1 2204 1 4 out_real_board_8[2]
rlabel metal3 3077 795 3077 795 4 out_real_board_8[1]
rlabel metal3 3077 1545 3077 1545 4 out_real_board_8[0]
rlabel metal3 3077 1595 3077 1595 4 out_real_board_9[2]
rlabel metal3 3077 1635 3077 1635 4 out_real_board_9[1]
rlabel metal3 3077 1485 3077 1485 4 out_real_board_9[0]
rlabel metal2 1708 3038 1708 3038 4 out_real_board_10[2]
rlabel metal2 1732 3038 1732 3038 4 out_real_board_10[1]
rlabel metal2 1692 3038 1692 3038 4 out_real_board_10[0]
rlabel metal3 3077 2325 3077 2325 4 out_real_board_11[2]
rlabel metal3 3077 2415 3077 2415 4 out_real_board_11[1]
rlabel metal3 3077 2525 3077 2525 4 out_real_board_11[0]
rlabel metal2 1836 3038 1836 3038 4 out_real_board_12[2]
rlabel metal2 2084 3038 2084 3038 4 out_real_board_12[1]
rlabel metal2 2068 3038 2068 3038 4 out_real_board_12[0]
rlabel metal2 2164 3038 2164 3038 4 out_real_board_13[2]
rlabel metal2 2324 3038 2324 3038 4 out_real_board_13[1]
rlabel metal3 3077 2305 3077 2305 4 out_real_board_13[0]
rlabel metal3 3077 1815 3077 1815 4 out_real_board_14[2]
rlabel metal3 3077 1725 3077 1725 4 out_real_board_14[1]
rlabel metal3 3077 1925 3077 1925 4 out_real_board_14[0]
rlabel metal3 3077 2125 3077 2125 4 out_real_board_15[2]
rlabel metal3 3077 1795 3077 1795 4 out_real_board_15[1]
rlabel metal3 3077 1615 3077 1615 4 out_real_board_15[0]
rlabel metal2 38 37 38 37 4 gnd
rlabel metal2 14 13 14 13 4 vdd
<< properties >>
string path 10404.000 26311.502 10404.000 26415.002 
<< end >>
